
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  n2491_lo,
  n2599_lo,
  n2611_lo,
  n2623_lo,
  n2635_lo,
  n2647_lo,
  n2659_lo,
  n2671_lo,
  n2683_lo,
  n2734_lo,
  n2746_lo,
  n2758_lo,
  n2770_lo,
  n2782_lo,
  n2794_lo,
  n2797_lo,
  n2806_lo,
  n2809_lo,
  n2818_lo,
  n2821_lo,
  n2830_lo,
  n2833_lo,
  n2839_lo,
  n2842_lo,
  n2845_lo,
  n2848_lo,
  n2851_lo,
  n2854_lo,
  n2857_lo,
  n2860_lo,
  n2863_lo,
  n3737_o2,
  n3736_o2,
  n3801_o2,
  n3836_o2,
  n3885_o2,
  n3902_o2,
  n4002_o2,
  n4052_o2,
  n4067_o2,
  n4162_o2,
  n4212_o2,
  n4227_o2,
  n4321_o2,
  n4367_o2,
  n4383_o2,
  n4475_o2,
  n4523_o2,
  n4537_o2,
  n4628_o2,
  n4674_o2,
  n4688_o2,
  n4791_o2,
  n4835_o2,
  n4868_o2,
  n5086_o2,
  n5130_o2,
  n5188_o2,
  n5402_o2,
  n5445_o2,
  n5500_o2,
  n5707_o2,
  n5745_o2,
  n5801_o2,
  n4836_o2,
  n4837_o2,
  n4838_o2,
  n4839_o2,
  n4840_o2,
  n4841_o2,
  n4842_o2,
  n4843_o2,
  n4844_o2,
  n4845_o2,
  n4846_o2,
  n4847_o2,
  n4848_o2,
  n4849_o2,
  n4850_o2,
  n4867_o2,
  n4908_o2,
  n6081_o2,
  n6120_o2,
  n316_inv,
  n4960_o2,
  n6203_o2,
  n325_inv,
  n328_inv,
  n331_inv,
  n5189_o2,
  n6594_o2,
  n340_inv,
  n6631_o2,
  n346_inv,
  n5388_o2,
  n6725_o2,
  n355_inv,
  n358_inv,
  n5612_o2,
  n1127_o2,
  n367_inv,
  n1231_o2,
  n373_inv,
  n5802_o2,
  n1232_o2,
  n382_inv,
  n385_inv,
  n6023_o2,
  n1235_o2,
  n394_inv,
  n1347_o2,
  n400_inv,
  n6383_o2,
  n1348_o2,
  n409_inv,
  n1351_o2,
  n1461_o2,
  n418_inv,
  n6024_o2,
  n6025_o2,
  n6026_o2,
  n6027_o2,
  n6028_o2,
  n6029_o2,
  n6030_o2,
  n6031_o2,
  n6032_o2,
  n6033_o2,
  n6034_o2,
  n6035_o2,
  n6036_o2,
  n6037_o2,
  n6038_o2,
  n6053_o2,
  n6726_o2,
  n6148_o2,
  n1463_o2,
  n1573_o2,
  n481_inv,
  n6201_o2,
  n487_inv,
  n490_inv,
  n493_inv,
  n1574_o2,
  n499_inv,
  n502_inv,
  n772_o2,
  n6482_o2,
  lo106_buf_o2,
  n1577_o2,
  n1678_o2,
  n520_inv,
  n523_inv,
  n6727_o2,
  n529_inv,
  n1679_o2,
  n535_inv,
  n848_o2,
  n541_inv,
  n544_inv,
  lo110_buf_o2,
  n1682_o2,
  n1775_o2,
  n512_o2,
  n559_inv,
  n562_inv,
  n2210_o2,
  n2126_o2,
  n2010_o2,
  n1776_o2,
  n577_inv,
  n580_inv,
  n932_o2,
  n548_o2,
  lo114_buf_o2,
  n1779_o2,
  n1864_o2,
  n598_inv,
  n601_inv,
  n592_o2,
  lo010_buf_o2,
  lo014_buf_o2,
  lo018_buf_o2,
  lo022_buf_o2,
  lo026_buf_o2,
  lo030_buf_o2,
  lo034_buf_o2,
  lo038_buf_o2,
  lo042_buf_o2,
  lo046_buf_o2,
  lo050_buf_o2,
  lo054_buf_o2,
  lo058_buf_o2,
  lo062_buf_o2,
  lo066_buf_o2,
  lo006_buf_o2,
  n655_inv,
  n2013_o2,
  n2129_o2,
  n2213_o2,
  n2243_o2,
  n2175_o2,
  n2075_o2,
  n1943_o2,
  n1865_o2,
  n682_inv,
  lo094_buf_o2,
  lo002_buf_o2,
  n691_inv,
  n451_o2,
  n1024_o2,
  n700_inv,
  n703_inv,
  n706_inv,
  lo118_buf_o2,
  n1868_o2,
  n1945_o2,
  n718_inv,
  n2045_o2,
  n1913_o2,
  n1749_o2,
  n1553_o2,
  n644_o2,
  n736_inv,
  lo098_buf_o2,
  n1121_o2,
  n1719_o2,
  n1523_o2,
  n464_o2,
  n754_inv,
  n757_inv,
  n760_inv,
  n2078_o2,
  n2079_o2,
  n2178_o2,
  n2179_o2,
  n2246_o2,
  n2247_o2,
  n2216_o2,
  n2217_o2,
  n2132_o2,
  n2133_o2,
  n2016_o2,
  n2017_o2,
  n1946_o2,
  n1556_o2,
  n1752_o2,
  n1916_o2,
  n2048_o2,
  n2102_o2,
  n1226_o2,
  n1986_o2,
  n1838_o2,
  n1658_o2,
  n829_inv,
  n1526_o2,
  n1722_o2,
  n1808_o2,
  n1628_o2,
  n844_inv,
  n847_inv,
  n1583_o2,
  n1787_o2,
  n1959_o2,
  n2099_o2,
  n2033_o2,
  n1877_o2,
  n1689_o2,
  n1355_o2,
  n1469_o2,
  n1238_o2,
  n1227_o2,
  n1124_o2,
  n704_o2,
  n484_o2,
  n1338_o2,
  n1449_o2,
  n1558_o2,
  n1754_o2,
  n1918_o2,
  n2050_o2,
  n2104_o2,
  n1988_o2,
  n1840_o2,
  n1660_o2,
  n708_o2,
  n768_o2,
  lo102_buf_o2,
  n1631_o2,
  n1632_o2,
  n1811_o2,
  n1812_o2,
  n1889_o2,
  n1890_o2,
  n1725_o2,
  n1726_o2,
  n917_o2,
  n918_o2,
  n1003_o2,
  n1004_o2,
  n1097_o2,
  n1098_o2,
  n1199_o2,
  n1200_o2,
  n1309_o2,
  n1310_o2,
  n1420_o2,
  n1421_o2,
  n1529_o2,
  n1530_o2,
  n839_o2,
  n840_o2,
  n577_o2,
  n623_o2,
  n677_o2,
  n739_o2,
  n809_o2,
  n887_o2,
  n973_o2,
  n1067_o2,
  n1169_o2,
  n1279_o2,
  n1390_o2,
  n1499_o2,
  n539_o2,
  lo082_buf_o2,
  n555_o2,
  n601_o2,
  n655_o2,
  n717_o2,
  n787_o2,
  n865_o2,
  n951_o2,
  n1045_o2,
  n1147_o2,
  n1257_o2,
  n1374_o2,
  n1488_o2,
  n1602_o2,
  n517_o2,
  n1603_o2,
  n509_o2,
  n510_o2,
  n579_o2,
  n625_o2,
  n679_o2,
  n741_o2,
  n811_o2,
  n889_o2,
  n975_o2,
  n1069_o2,
  n1171_o2,
  n1281_o2,
  n1392_o2,
  n1501_o2,
  n541_o2,
  G6257,
  G6258,
  G6259,
  G6260,
  G6261,
  G6262,
  G6263,
  G6264,
  G6265,
  G6266,
  G6267,
  G6268,
  G6269,
  G6270,
  G6271,
  G6272,
  G6273,
  G6274,
  G6275,
  G6276,
  G6277,
  G6278,
  G6279,
  G6280,
  G6281,
  G6282,
  G6283,
  G6284,
  G6285,
  G6286,
  G6287,
  G6288,
  n5322_li003_li003,
  n5430_li039_li039,
  n5442_li043_li043,
  n5454_li047_li047,
  n5466_li051_li051,
  n5478_li055_li055,
  n5490_li059_li059,
  n5502_li063_li063,
  n5514_li067_li067,
  n5565_li084_li084,
  n5577_li088_li088,
  n5589_li092_li092,
  n5601_li096_li096,
  n5613_li100_li100,
  n5625_li104_li104,
  n5628_li105_li105,
  n5637_li108_li108,
  n5640_li109_li109,
  n5649_li112_li112,
  n5652_li113_li113,
  n5661_li116_li116,
  n5664_li117_li117,
  n5670_li119_li119,
  n5673_li120_li120,
  n5676_li121_li121,
  n5679_li122_li122,
  n5682_li123_li123,
  n5685_li124_li124,
  n5688_li125_li125,
  n5691_li126_li126,
  n5694_li127_li127,
  n3737_i2,
  n3736_i2,
  n3801_i2,
  n3836_i2,
  n3885_i2,
  n3902_i2,
  n4002_i2,
  n4052_i2,
  n4067_i2,
  n4162_i2,
  n4212_i2,
  n4227_i2,
  n4321_i2,
  n4367_i2,
  n4383_i2,
  n4475_i2,
  n4523_i2,
  n4537_i2,
  n4628_i2,
  n4674_i2,
  n4688_i2,
  n4791_i2,
  n4835_i2,
  n4868_i2,
  n5086_i2,
  n5130_i2,
  n5188_i2,
  n5402_i2,
  n5445_i2,
  n5500_i2,
  n5707_i2,
  n5745_i2,
  n5801_i2,
  n4836_i2,
  n4837_i2,
  n4838_i2,
  n4839_i2,
  n4840_i2,
  n4841_i2,
  n4842_i2,
  n4843_i2,
  n4844_i2,
  n4845_i2,
  n4846_i2,
  n4847_i2,
  n4848_i2,
  n4849_i2,
  n4850_i2,
  n4867_i2,
  n4908_i2,
  n6081_i2,
  n6120_i2,
  n4959_i2,
  n4960_i2,
  n6203_i2,
  n5040_i2,
  n5087_i2,
  n5158_i2,
  n5189_i2,
  n6594_i2,
  n5328_i2,
  n6631_i2,
  n5372_i2,
  n5388_i2,
  n6725_i2,
  n5527_i2,
  n5555_i2,
  n5612_i2,
  n1127_i2,
  n5708_i2,
  n1231_i2,
  n5771_i2,
  n5802_i2,
  n1232_i2,
  n5948_i2,
  n6006_i2,
  n6023_i2,
  n1235_i2,
  n6243_i2,
  n1347_i2,
  n6296_i2,
  n6383_i2,
  n1348_i2,
  n6595_i2,
  n1351_i2,
  n1461_i2,
  n6655_i2,
  n6024_i2,
  n6025_i2,
  n6026_i2,
  n6027_i2,
  n6028_i2,
  n6029_i2,
  n6030_i2,
  n6031_i2,
  n6032_i2,
  n6033_i2,
  n6034_i2,
  n6035_i2,
  n6036_i2,
  n6037_i2,
  n6038_i2,
  n6053_i2,
  n6726_i2,
  n6148_i2,
  n1463_i2,
  n1573_i2,
  n6200_i2,
  n6201_i2,
  n6294_i2,
  n707_i2,
  n6361_i2,
  n1574_i2,
  n771_i2,
  n6423_i2,
  n772_i2,
  n6482_i2,
  lo106_buf_i2,
  n1577_i2,
  n1678_i2,
  n6596_i2,
  n6683_i2,
  n6727_i2,
  n775_i2,
  n1679_i2,
  n847_i2,
  n848_i2,
  n487_i2,
  n511_i2,
  lo110_buf_i2,
  n1682_i2,
  n1775_i2,
  n512_i2,
  n851_i2,
  n515_i2,
  n2210_i2,
  n2126_i2,
  n2010_i2,
  n1776_i2,
  n931_i2,
  n547_i2,
  n932_i2,
  n548_i2,
  lo114_buf_i2,
  n1779_i2,
  n1864_i2,
  n551_i2,
  n591_i2,
  n592_i2,
  lo010_buf_i2,
  lo014_buf_i2,
  lo018_buf_i2,
  lo022_buf_i2,
  lo026_buf_i2,
  lo030_buf_i2,
  lo034_buf_i2,
  lo038_buf_i2,
  lo042_buf_i2,
  lo046_buf_i2,
  lo050_buf_i2,
  lo054_buf_i2,
  lo058_buf_i2,
  lo062_buf_i2,
  lo066_buf_i2,
  lo006_buf_i2,
  n935_i2,
  n2013_i2,
  n2129_i2,
  n2213_i2,
  n2243_i2,
  n2175_i2,
  n2075_i2,
  n1943_i2,
  n1865_i2,
  n1023_i2,
  lo094_buf_i2,
  lo002_buf_i2,
  n450_i2,
  n451_i2,
  n1024_i2,
  n595_i2,
  n452_i2,
  n643_i2,
  lo118_buf_i2,
  n1868_i2,
  n1945_i2,
  n455_i2,
  n2045_i2,
  n1913_i2,
  n1749_i2,
  n1553_i2,
  n644_i2,
  n463_i2,
  lo098_buf_i2,
  n1121_i2,
  n1719_i2,
  n1523_i2,
  n464_i2,
  n1027_i2,
  n647_i2,
  n467_i2,
  n2078_i2,
  n2079_i2,
  n2178_i2,
  n2179_i2,
  n2246_i2,
  n2247_i2,
  n2216_i2,
  n2217_i2,
  n2132_i2,
  n2133_i2,
  n2016_i2,
  n2017_i2,
  n1946_i2,
  n1556_i2,
  n1752_i2,
  n1916_i2,
  n2048_i2,
  n2102_i2,
  n1226_i2,
  n1986_i2,
  n1838_i2,
  n1658_i2,
  n1123_i2,
  n1526_i2,
  n1722_i2,
  n1808_i2,
  n1628_i2,
  n703_i2,
  n483_i2,
  n1583_i2,
  n1787_i2,
  n1959_i2,
  n2099_i2,
  n2033_i2,
  n1877_i2,
  n1689_i2,
  n1355_i2,
  n1469_i2,
  n1238_i2,
  n1227_i2,
  n1124_i2,
  n704_i2,
  n484_i2,
  n1338_i2,
  n1449_i2,
  n1558_i2,
  n1754_i2,
  n1918_i2,
  n2050_i2,
  n2104_i2,
  n1988_i2,
  n1840_i2,
  n1660_i2,
  n708_i2,
  n768_i2,
  lo102_buf_i2,
  n1631_i2,
  n1632_i2,
  n1811_i2,
  n1812_i2,
  n1889_i2,
  n1890_i2,
  n1725_i2,
  n1726_i2,
  n917_i2,
  n918_i2,
  n1003_i2,
  n1004_i2,
  n1097_i2,
  n1098_i2,
  n1199_i2,
  n1200_i2,
  n1309_i2,
  n1310_i2,
  n1420_i2,
  n1421_i2,
  n1529_i2,
  n1530_i2,
  n839_i2,
  n840_i2,
  n577_i2,
  n623_i2,
  n677_i2,
  n739_i2,
  n809_i2,
  n887_i2,
  n973_i2,
  n1067_i2,
  n1169_i2,
  n1279_i2,
  n1390_i2,
  n1499_i2,
  n539_i2,
  lo082_buf_i2,
  n555_i2,
  n601_i2,
  n655_i2,
  n717_i2,
  n787_i2,
  n865_i2,
  n951_i2,
  n1045_i2,
  n1147_i2,
  n1257_i2,
  n1374_i2,
  n1488_i2,
  n1602_i2,
  n517_i2,
  n1603_i2,
  n509_i2,
  n510_i2,
  n579_i2,
  n625_i2,
  n679_i2,
  n741_i2,
  n811_i2,
  n889_i2,
  n975_i2,
  n1069_i2,
  n1171_i2,
  n1281_i2,
  n1392_i2,
  n1501_i2,
  n541_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input n2491_lo;input n2599_lo;input n2611_lo;input n2623_lo;input n2635_lo;input n2647_lo;input n2659_lo;input n2671_lo;input n2683_lo;input n2734_lo;input n2746_lo;input n2758_lo;input n2770_lo;input n2782_lo;input n2794_lo;input n2797_lo;input n2806_lo;input n2809_lo;input n2818_lo;input n2821_lo;input n2830_lo;input n2833_lo;input n2839_lo;input n2842_lo;input n2845_lo;input n2848_lo;input n2851_lo;input n2854_lo;input n2857_lo;input n2860_lo;input n2863_lo;input n3737_o2;input n3736_o2;input n3801_o2;input n3836_o2;input n3885_o2;input n3902_o2;input n4002_o2;input n4052_o2;input n4067_o2;input n4162_o2;input n4212_o2;input n4227_o2;input n4321_o2;input n4367_o2;input n4383_o2;input n4475_o2;input n4523_o2;input n4537_o2;input n4628_o2;input n4674_o2;input n4688_o2;input n4791_o2;input n4835_o2;input n4868_o2;input n5086_o2;input n5130_o2;input n5188_o2;input n5402_o2;input n5445_o2;input n5500_o2;input n5707_o2;input n5745_o2;input n5801_o2;input n4836_o2;input n4837_o2;input n4838_o2;input n4839_o2;input n4840_o2;input n4841_o2;input n4842_o2;input n4843_o2;input n4844_o2;input n4845_o2;input n4846_o2;input n4847_o2;input n4848_o2;input n4849_o2;input n4850_o2;input n4867_o2;input n4908_o2;input n6081_o2;input n6120_o2;input n316_inv;input n4960_o2;input n6203_o2;input n325_inv;input n328_inv;input n331_inv;input n5189_o2;input n6594_o2;input n340_inv;input n6631_o2;input n346_inv;input n5388_o2;input n6725_o2;input n355_inv;input n358_inv;input n5612_o2;input n1127_o2;input n367_inv;input n1231_o2;input n373_inv;input n5802_o2;input n1232_o2;input n382_inv;input n385_inv;input n6023_o2;input n1235_o2;input n394_inv;input n1347_o2;input n400_inv;input n6383_o2;input n1348_o2;input n409_inv;input n1351_o2;input n1461_o2;input n418_inv;input n6024_o2;input n6025_o2;input n6026_o2;input n6027_o2;input n6028_o2;input n6029_o2;input n6030_o2;input n6031_o2;input n6032_o2;input n6033_o2;input n6034_o2;input n6035_o2;input n6036_o2;input n6037_o2;input n6038_o2;input n6053_o2;input n6726_o2;input n6148_o2;input n1463_o2;input n1573_o2;input n481_inv;input n6201_o2;input n487_inv;input n490_inv;input n493_inv;input n1574_o2;input n499_inv;input n502_inv;input n772_o2;input n6482_o2;input lo106_buf_o2;input n1577_o2;input n1678_o2;input n520_inv;input n523_inv;input n6727_o2;input n529_inv;input n1679_o2;input n535_inv;input n848_o2;input n541_inv;input n544_inv;input lo110_buf_o2;input n1682_o2;input n1775_o2;input n512_o2;input n559_inv;input n562_inv;input n2210_o2;input n2126_o2;input n2010_o2;input n1776_o2;input n577_inv;input n580_inv;input n932_o2;input n548_o2;input lo114_buf_o2;input n1779_o2;input n1864_o2;input n598_inv;input n601_inv;input n592_o2;input lo010_buf_o2;input lo014_buf_o2;input lo018_buf_o2;input lo022_buf_o2;input lo026_buf_o2;input lo030_buf_o2;input lo034_buf_o2;input lo038_buf_o2;input lo042_buf_o2;input lo046_buf_o2;input lo050_buf_o2;input lo054_buf_o2;input lo058_buf_o2;input lo062_buf_o2;input lo066_buf_o2;input lo006_buf_o2;input n655_inv;input n2013_o2;input n2129_o2;input n2213_o2;input n2243_o2;input n2175_o2;input n2075_o2;input n1943_o2;input n1865_o2;input n682_inv;input lo094_buf_o2;input lo002_buf_o2;input n691_inv;input n451_o2;input n1024_o2;input n700_inv;input n703_inv;input n706_inv;input lo118_buf_o2;input n1868_o2;input n1945_o2;input n718_inv;input n2045_o2;input n1913_o2;input n1749_o2;input n1553_o2;input n644_o2;input n736_inv;input lo098_buf_o2;input n1121_o2;input n1719_o2;input n1523_o2;input n464_o2;input n754_inv;input n757_inv;input n760_inv;input n2078_o2;input n2079_o2;input n2178_o2;input n2179_o2;input n2246_o2;input n2247_o2;input n2216_o2;input n2217_o2;input n2132_o2;input n2133_o2;input n2016_o2;input n2017_o2;input n1946_o2;input n1556_o2;input n1752_o2;input n1916_o2;input n2048_o2;input n2102_o2;input n1226_o2;input n1986_o2;input n1838_o2;input n1658_o2;input n829_inv;input n1526_o2;input n1722_o2;input n1808_o2;input n1628_o2;input n844_inv;input n847_inv;input n1583_o2;input n1787_o2;input n1959_o2;input n2099_o2;input n2033_o2;input n1877_o2;input n1689_o2;input n1355_o2;input n1469_o2;input n1238_o2;input n1227_o2;input n1124_o2;input n704_o2;input n484_o2;input n1338_o2;input n1449_o2;input n1558_o2;input n1754_o2;input n1918_o2;input n2050_o2;input n2104_o2;input n1988_o2;input n1840_o2;input n1660_o2;input n708_o2;input n768_o2;input lo102_buf_o2;input n1631_o2;input n1632_o2;input n1811_o2;input n1812_o2;input n1889_o2;input n1890_o2;input n1725_o2;input n1726_o2;input n917_o2;input n918_o2;input n1003_o2;input n1004_o2;input n1097_o2;input n1098_o2;input n1199_o2;input n1200_o2;input n1309_o2;input n1310_o2;input n1420_o2;input n1421_o2;input n1529_o2;input n1530_o2;input n839_o2;input n840_o2;input n577_o2;input n623_o2;input n677_o2;input n739_o2;input n809_o2;input n887_o2;input n973_o2;input n1067_o2;input n1169_o2;input n1279_o2;input n1390_o2;input n1499_o2;input n539_o2;input lo082_buf_o2;input n555_o2;input n601_o2;input n655_o2;input n717_o2;input n787_o2;input n865_o2;input n951_o2;input n1045_o2;input n1147_o2;input n1257_o2;input n1374_o2;input n1488_o2;input n1602_o2;input n517_o2;input n1603_o2;input n509_o2;input n510_o2;input n579_o2;input n625_o2;input n679_o2;input n741_o2;input n811_o2;input n889_o2;input n975_o2;input n1069_o2;input n1171_o2;input n1281_o2;input n1392_o2;input n1501_o2;input n541_o2;
  output G6257;output G6258;output G6259;output G6260;output G6261;output G6262;output G6263;output G6264;output G6265;output G6266;output G6267;output G6268;output G6269;output G6270;output G6271;output G6272;output G6273;output G6274;output G6275;output G6276;output G6277;output G6278;output G6279;output G6280;output G6281;output G6282;output G6283;output G6284;output G6285;output G6286;output G6287;output G6288;output n5322_li003_li003;output n5430_li039_li039;output n5442_li043_li043;output n5454_li047_li047;output n5466_li051_li051;output n5478_li055_li055;output n5490_li059_li059;output n5502_li063_li063;output n5514_li067_li067;output n5565_li084_li084;output n5577_li088_li088;output n5589_li092_li092;output n5601_li096_li096;output n5613_li100_li100;output n5625_li104_li104;output n5628_li105_li105;output n5637_li108_li108;output n5640_li109_li109;output n5649_li112_li112;output n5652_li113_li113;output n5661_li116_li116;output n5664_li117_li117;output n5670_li119_li119;output n5673_li120_li120;output n5676_li121_li121;output n5679_li122_li122;output n5682_li123_li123;output n5685_li124_li124;output n5688_li125_li125;output n5691_li126_li126;output n5694_li127_li127;output n3737_i2;output n3736_i2;output n3801_i2;output n3836_i2;output n3885_i2;output n3902_i2;output n4002_i2;output n4052_i2;output n4067_i2;output n4162_i2;output n4212_i2;output n4227_i2;output n4321_i2;output n4367_i2;output n4383_i2;output n4475_i2;output n4523_i2;output n4537_i2;output n4628_i2;output n4674_i2;output n4688_i2;output n4791_i2;output n4835_i2;output n4868_i2;output n5086_i2;output n5130_i2;output n5188_i2;output n5402_i2;output n5445_i2;output n5500_i2;output n5707_i2;output n5745_i2;output n5801_i2;output n4836_i2;output n4837_i2;output n4838_i2;output n4839_i2;output n4840_i2;output n4841_i2;output n4842_i2;output n4843_i2;output n4844_i2;output n4845_i2;output n4846_i2;output n4847_i2;output n4848_i2;output n4849_i2;output n4850_i2;output n4867_i2;output n4908_i2;output n6081_i2;output n6120_i2;output n4959_i2;output n4960_i2;output n6203_i2;output n5040_i2;output n5087_i2;output n5158_i2;output n5189_i2;output n6594_i2;output n5328_i2;output n6631_i2;output n5372_i2;output n5388_i2;output n6725_i2;output n5527_i2;output n5555_i2;output n5612_i2;output n1127_i2;output n5708_i2;output n1231_i2;output n5771_i2;output n5802_i2;output n1232_i2;output n5948_i2;output n6006_i2;output n6023_i2;output n1235_i2;output n6243_i2;output n1347_i2;output n6296_i2;output n6383_i2;output n1348_i2;output n6595_i2;output n1351_i2;output n1461_i2;output n6655_i2;output n6024_i2;output n6025_i2;output n6026_i2;output n6027_i2;output n6028_i2;output n6029_i2;output n6030_i2;output n6031_i2;output n6032_i2;output n6033_i2;output n6034_i2;output n6035_i2;output n6036_i2;output n6037_i2;output n6038_i2;output n6053_i2;output n6726_i2;output n6148_i2;output n1463_i2;output n1573_i2;output n6200_i2;output n6201_i2;output n6294_i2;output n707_i2;output n6361_i2;output n1574_i2;output n771_i2;output n6423_i2;output n772_i2;output n6482_i2;output lo106_buf_i2;output n1577_i2;output n1678_i2;output n6596_i2;output n6683_i2;output n6727_i2;output n775_i2;output n1679_i2;output n847_i2;output n848_i2;output n487_i2;output n511_i2;output lo110_buf_i2;output n1682_i2;output n1775_i2;output n512_i2;output n851_i2;output n515_i2;output n2210_i2;output n2126_i2;output n2010_i2;output n1776_i2;output n931_i2;output n547_i2;output n932_i2;output n548_i2;output lo114_buf_i2;output n1779_i2;output n1864_i2;output n551_i2;output n591_i2;output n592_i2;output lo010_buf_i2;output lo014_buf_i2;output lo018_buf_i2;output lo022_buf_i2;output lo026_buf_i2;output lo030_buf_i2;output lo034_buf_i2;output lo038_buf_i2;output lo042_buf_i2;output lo046_buf_i2;output lo050_buf_i2;output lo054_buf_i2;output lo058_buf_i2;output lo062_buf_i2;output lo066_buf_i2;output lo006_buf_i2;output n935_i2;output n2013_i2;output n2129_i2;output n2213_i2;output n2243_i2;output n2175_i2;output n2075_i2;output n1943_i2;output n1865_i2;output n1023_i2;output lo094_buf_i2;output lo002_buf_i2;output n450_i2;output n451_i2;output n1024_i2;output n595_i2;output n452_i2;output n643_i2;output lo118_buf_i2;output n1868_i2;output n1945_i2;output n455_i2;output n2045_i2;output n1913_i2;output n1749_i2;output n1553_i2;output n644_i2;output n463_i2;output lo098_buf_i2;output n1121_i2;output n1719_i2;output n1523_i2;output n464_i2;output n1027_i2;output n647_i2;output n467_i2;output n2078_i2;output n2079_i2;output n2178_i2;output n2179_i2;output n2246_i2;output n2247_i2;output n2216_i2;output n2217_i2;output n2132_i2;output n2133_i2;output n2016_i2;output n2017_i2;output n1946_i2;output n1556_i2;output n1752_i2;output n1916_i2;output n2048_i2;output n2102_i2;output n1226_i2;output n1986_i2;output n1838_i2;output n1658_i2;output n1123_i2;output n1526_i2;output n1722_i2;output n1808_i2;output n1628_i2;output n703_i2;output n483_i2;output n1583_i2;output n1787_i2;output n1959_i2;output n2099_i2;output n2033_i2;output n1877_i2;output n1689_i2;output n1355_i2;output n1469_i2;output n1238_i2;output n1227_i2;output n1124_i2;output n704_i2;output n484_i2;output n1338_i2;output n1449_i2;output n1558_i2;output n1754_i2;output n1918_i2;output n2050_i2;output n2104_i2;output n1988_i2;output n1840_i2;output n1660_i2;output n708_i2;output n768_i2;output lo102_buf_i2;output n1631_i2;output n1632_i2;output n1811_i2;output n1812_i2;output n1889_i2;output n1890_i2;output n1725_i2;output n1726_i2;output n917_i2;output n918_i2;output n1003_i2;output n1004_i2;output n1097_i2;output n1098_i2;output n1199_i2;output n1200_i2;output n1309_i2;output n1310_i2;output n1420_i2;output n1421_i2;output n1529_i2;output n1530_i2;output n839_i2;output n840_i2;output n577_i2;output n623_i2;output n677_i2;output n739_i2;output n809_i2;output n887_i2;output n973_i2;output n1067_i2;output n1169_i2;output n1279_i2;output n1390_i2;output n1499_i2;output n539_i2;output lo082_buf_i2;output n555_i2;output n601_i2;output n655_i2;output n717_i2;output n787_i2;output n865_i2;output n951_i2;output n1045_i2;output n1147_i2;output n1257_i2;output n1374_i2;output n1488_i2;output n1602_i2;output n517_i2;output n1603_i2;output n509_i2;output n510_i2;output n579_i2;output n625_i2;output n679_i2;output n741_i2;output n811_i2;output n889_i2;output n975_i2;output n1069_i2;output n1171_i2;output n1281_i2;output n1392_i2;output n1501_i2;output n541_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire n2491_lo_p;
  wire n2491_lo_n;
  wire n2599_lo_p;
  wire n2599_lo_n;
  wire n2611_lo_p;
  wire n2611_lo_n;
  wire n2623_lo_p;
  wire n2623_lo_n;
  wire n2635_lo_p;
  wire n2635_lo_n;
  wire n2647_lo_p;
  wire n2647_lo_n;
  wire n2659_lo_p;
  wire n2659_lo_n;
  wire n2671_lo_p;
  wire n2671_lo_n;
  wire n2683_lo_p;
  wire n2683_lo_n;
  wire n2734_lo_p;
  wire n2734_lo_n;
  wire n2746_lo_p;
  wire n2746_lo_n;
  wire n2758_lo_p;
  wire n2758_lo_n;
  wire n2770_lo_p;
  wire n2770_lo_n;
  wire n2782_lo_p;
  wire n2782_lo_n;
  wire n2794_lo_p;
  wire n2794_lo_n;
  wire n2797_lo_p;
  wire n2797_lo_n;
  wire n2806_lo_p;
  wire n2806_lo_n;
  wire n2809_lo_p;
  wire n2809_lo_n;
  wire n2818_lo_p;
  wire n2818_lo_n;
  wire n2821_lo_p;
  wire n2821_lo_n;
  wire n2830_lo_p;
  wire n2830_lo_n;
  wire n2833_lo_p;
  wire n2833_lo_n;
  wire n2839_lo_p;
  wire n2839_lo_n;
  wire n2842_lo_p;
  wire n2842_lo_n;
  wire n2845_lo_p;
  wire n2845_lo_n;
  wire n2848_lo_p;
  wire n2848_lo_n;
  wire n2851_lo_p;
  wire n2851_lo_n;
  wire n2854_lo_p;
  wire n2854_lo_n;
  wire n2857_lo_p;
  wire n2857_lo_n;
  wire n2860_lo_p;
  wire n2860_lo_n;
  wire n2863_lo_p;
  wire n2863_lo_n;
  wire n3737_o2_p;
  wire n3737_o2_n;
  wire n3736_o2_p;
  wire n3736_o2_n;
  wire n3801_o2_p;
  wire n3801_o2_n;
  wire n3836_o2_p;
  wire n3836_o2_n;
  wire n3885_o2_p;
  wire n3885_o2_n;
  wire n3902_o2_p;
  wire n3902_o2_n;
  wire n4002_o2_p;
  wire n4002_o2_n;
  wire n4052_o2_p;
  wire n4052_o2_n;
  wire n4067_o2_p;
  wire n4067_o2_n;
  wire n4162_o2_p;
  wire n4162_o2_n;
  wire n4212_o2_p;
  wire n4212_o2_n;
  wire n4227_o2_p;
  wire n4227_o2_n;
  wire n4321_o2_p;
  wire n4321_o2_n;
  wire n4367_o2_p;
  wire n4367_o2_n;
  wire n4383_o2_p;
  wire n4383_o2_n;
  wire n4475_o2_p;
  wire n4475_o2_n;
  wire n4523_o2_p;
  wire n4523_o2_n;
  wire n4537_o2_p;
  wire n4537_o2_n;
  wire n4628_o2_p;
  wire n4628_o2_n;
  wire n4674_o2_p;
  wire n4674_o2_n;
  wire n4688_o2_p;
  wire n4688_o2_n;
  wire n4791_o2_p;
  wire n4791_o2_n;
  wire n4835_o2_p;
  wire n4835_o2_n;
  wire n4868_o2_p;
  wire n4868_o2_n;
  wire n5086_o2_p;
  wire n5086_o2_n;
  wire n5130_o2_p;
  wire n5130_o2_n;
  wire n5188_o2_p;
  wire n5188_o2_n;
  wire n5402_o2_p;
  wire n5402_o2_n;
  wire n5445_o2_p;
  wire n5445_o2_n;
  wire n5500_o2_p;
  wire n5500_o2_n;
  wire n5707_o2_p;
  wire n5707_o2_n;
  wire n5745_o2_p;
  wire n5745_o2_n;
  wire n5801_o2_p;
  wire n5801_o2_n;
  wire n4836_o2_p;
  wire n4836_o2_n;
  wire n4837_o2_p;
  wire n4837_o2_n;
  wire n4838_o2_p;
  wire n4838_o2_n;
  wire n4839_o2_p;
  wire n4839_o2_n;
  wire n4840_o2_p;
  wire n4840_o2_n;
  wire n4841_o2_p;
  wire n4841_o2_n;
  wire n4842_o2_p;
  wire n4842_o2_n;
  wire n4843_o2_p;
  wire n4843_o2_n;
  wire n4844_o2_p;
  wire n4844_o2_n;
  wire n4845_o2_p;
  wire n4845_o2_n;
  wire n4846_o2_p;
  wire n4846_o2_n;
  wire n4847_o2_p;
  wire n4847_o2_n;
  wire n4848_o2_p;
  wire n4848_o2_n;
  wire n4849_o2_p;
  wire n4849_o2_n;
  wire n4850_o2_p;
  wire n4850_o2_n;
  wire n4867_o2_p;
  wire n4867_o2_n;
  wire n4908_o2_p;
  wire n4908_o2_n;
  wire n6081_o2_p;
  wire n6081_o2_n;
  wire n6120_o2_p;
  wire n6120_o2_n;
  wire n316_inv_p;
  wire n316_inv_n;
  wire n4960_o2_p;
  wire n4960_o2_n;
  wire n6203_o2_p;
  wire n6203_o2_n;
  wire n325_inv_p;
  wire n325_inv_n;
  wire n328_inv_p;
  wire n328_inv_n;
  wire n331_inv_p;
  wire n331_inv_n;
  wire n5189_o2_p;
  wire n5189_o2_n;
  wire n6594_o2_p;
  wire n6594_o2_n;
  wire n340_inv_p;
  wire n340_inv_n;
  wire n6631_o2_p;
  wire n6631_o2_n;
  wire n346_inv_p;
  wire n346_inv_n;
  wire n5388_o2_p;
  wire n5388_o2_n;
  wire n6725_o2_p;
  wire n6725_o2_n;
  wire n355_inv_p;
  wire n355_inv_n;
  wire n358_inv_p;
  wire n358_inv_n;
  wire n5612_o2_p;
  wire n5612_o2_n;
  wire n1127_o2_p;
  wire n1127_o2_n;
  wire n367_inv_p;
  wire n367_inv_n;
  wire n1231_o2_p;
  wire n1231_o2_n;
  wire n373_inv_p;
  wire n373_inv_n;
  wire n5802_o2_p;
  wire n5802_o2_n;
  wire n1232_o2_p;
  wire n1232_o2_n;
  wire n382_inv_p;
  wire n382_inv_n;
  wire n385_inv_p;
  wire n385_inv_n;
  wire n6023_o2_p;
  wire n6023_o2_n;
  wire n1235_o2_p;
  wire n1235_o2_n;
  wire n394_inv_p;
  wire n394_inv_n;
  wire n1347_o2_p;
  wire n1347_o2_n;
  wire n400_inv_p;
  wire n400_inv_n;
  wire n6383_o2_p;
  wire n6383_o2_n;
  wire n1348_o2_p;
  wire n1348_o2_n;
  wire n409_inv_p;
  wire n409_inv_n;
  wire n1351_o2_p;
  wire n1351_o2_n;
  wire n1461_o2_p;
  wire n1461_o2_n;
  wire n418_inv_p;
  wire n418_inv_n;
  wire n6024_o2_p;
  wire n6024_o2_n;
  wire n6025_o2_p;
  wire n6025_o2_n;
  wire n6026_o2_p;
  wire n6026_o2_n;
  wire n6027_o2_p;
  wire n6027_o2_n;
  wire n6028_o2_p;
  wire n6028_o2_n;
  wire n6029_o2_p;
  wire n6029_o2_n;
  wire n6030_o2_p;
  wire n6030_o2_n;
  wire n6031_o2_p;
  wire n6031_o2_n;
  wire n6032_o2_p;
  wire n6032_o2_n;
  wire n6033_o2_p;
  wire n6033_o2_n;
  wire n6034_o2_p;
  wire n6034_o2_n;
  wire n6035_o2_p;
  wire n6035_o2_n;
  wire n6036_o2_p;
  wire n6036_o2_n;
  wire n6037_o2_p;
  wire n6037_o2_n;
  wire n6038_o2_p;
  wire n6038_o2_n;
  wire n6053_o2_p;
  wire n6053_o2_n;
  wire n6726_o2_p;
  wire n6726_o2_n;
  wire n6148_o2_p;
  wire n6148_o2_n;
  wire n1463_o2_p;
  wire n1463_o2_n;
  wire n1573_o2_p;
  wire n1573_o2_n;
  wire n481_inv_p;
  wire n481_inv_n;
  wire n6201_o2_p;
  wire n6201_o2_n;
  wire n487_inv_p;
  wire n487_inv_n;
  wire n490_inv_p;
  wire n490_inv_n;
  wire n493_inv_p;
  wire n493_inv_n;
  wire n1574_o2_p;
  wire n1574_o2_n;
  wire n499_inv_p;
  wire n499_inv_n;
  wire n502_inv_p;
  wire n502_inv_n;
  wire n772_o2_p;
  wire n772_o2_n;
  wire n6482_o2_p;
  wire n6482_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire n1577_o2_p;
  wire n1577_o2_n;
  wire n1678_o2_p;
  wire n1678_o2_n;
  wire n520_inv_p;
  wire n520_inv_n;
  wire n523_inv_p;
  wire n523_inv_n;
  wire n6727_o2_p;
  wire n6727_o2_n;
  wire n529_inv_p;
  wire n529_inv_n;
  wire n1679_o2_p;
  wire n1679_o2_n;
  wire n535_inv_p;
  wire n535_inv_n;
  wire n848_o2_p;
  wire n848_o2_n;
  wire n541_inv_p;
  wire n541_inv_n;
  wire n544_inv_p;
  wire n544_inv_n;
  wire lo110_buf_o2_p;
  wire lo110_buf_o2_n;
  wire n1682_o2_p;
  wire n1682_o2_n;
  wire n1775_o2_p;
  wire n1775_o2_n;
  wire n512_o2_p;
  wire n512_o2_n;
  wire n559_inv_p;
  wire n559_inv_n;
  wire n562_inv_p;
  wire n562_inv_n;
  wire n2210_o2_p;
  wire n2210_o2_n;
  wire n2126_o2_p;
  wire n2126_o2_n;
  wire n2010_o2_p;
  wire n2010_o2_n;
  wire n1776_o2_p;
  wire n1776_o2_n;
  wire n577_inv_p;
  wire n577_inv_n;
  wire n580_inv_p;
  wire n580_inv_n;
  wire n932_o2_p;
  wire n932_o2_n;
  wire n548_o2_p;
  wire n548_o2_n;
  wire lo114_buf_o2_p;
  wire lo114_buf_o2_n;
  wire n1779_o2_p;
  wire n1779_o2_n;
  wire n1864_o2_p;
  wire n1864_o2_n;
  wire n598_inv_p;
  wire n598_inv_n;
  wire n601_inv_p;
  wire n601_inv_n;
  wire n592_o2_p;
  wire n592_o2_n;
  wire lo010_buf_o2_p;
  wire lo010_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo018_buf_o2_p;
  wire lo018_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo026_buf_o2_p;
  wire lo026_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo034_buf_o2_p;
  wire lo034_buf_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo046_buf_o2_p;
  wire lo046_buf_o2_n;
  wire lo050_buf_o2_p;
  wire lo050_buf_o2_n;
  wire lo054_buf_o2_p;
  wire lo054_buf_o2_n;
  wire lo058_buf_o2_p;
  wire lo058_buf_o2_n;
  wire lo062_buf_o2_p;
  wire lo062_buf_o2_n;
  wire lo066_buf_o2_p;
  wire lo066_buf_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire n655_inv_p;
  wire n655_inv_n;
  wire n2013_o2_p;
  wire n2013_o2_n;
  wire n2129_o2_p;
  wire n2129_o2_n;
  wire n2213_o2_p;
  wire n2213_o2_n;
  wire n2243_o2_p;
  wire n2243_o2_n;
  wire n2175_o2_p;
  wire n2175_o2_n;
  wire n2075_o2_p;
  wire n2075_o2_n;
  wire n1943_o2_p;
  wire n1943_o2_n;
  wire n1865_o2_p;
  wire n1865_o2_n;
  wire n682_inv_p;
  wire n682_inv_n;
  wire lo094_buf_o2_p;
  wire lo094_buf_o2_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire n691_inv_p;
  wire n691_inv_n;
  wire n451_o2_p;
  wire n451_o2_n;
  wire n1024_o2_p;
  wire n1024_o2_n;
  wire n700_inv_p;
  wire n700_inv_n;
  wire n703_inv_p;
  wire n703_inv_n;
  wire n706_inv_p;
  wire n706_inv_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire n1868_o2_p;
  wire n1868_o2_n;
  wire n1945_o2_p;
  wire n1945_o2_n;
  wire n718_inv_p;
  wire n718_inv_n;
  wire n2045_o2_p;
  wire n2045_o2_n;
  wire n1913_o2_p;
  wire n1913_o2_n;
  wire n1749_o2_p;
  wire n1749_o2_n;
  wire n1553_o2_p;
  wire n1553_o2_n;
  wire n644_o2_p;
  wire n644_o2_n;
  wire n736_inv_p;
  wire n736_inv_n;
  wire lo098_buf_o2_p;
  wire lo098_buf_o2_n;
  wire n1121_o2_p;
  wire n1121_o2_n;
  wire n1719_o2_p;
  wire n1719_o2_n;
  wire n1523_o2_p;
  wire n1523_o2_n;
  wire n464_o2_p;
  wire n464_o2_n;
  wire n754_inv_p;
  wire n754_inv_n;
  wire n757_inv_p;
  wire n757_inv_n;
  wire n760_inv_p;
  wire n760_inv_n;
  wire n2078_o2_p;
  wire n2078_o2_n;
  wire n2079_o2_p;
  wire n2079_o2_n;
  wire n2178_o2_p;
  wire n2178_o2_n;
  wire n2179_o2_p;
  wire n2179_o2_n;
  wire n2246_o2_p;
  wire n2246_o2_n;
  wire n2247_o2_p;
  wire n2247_o2_n;
  wire n2216_o2_p;
  wire n2216_o2_n;
  wire n2217_o2_p;
  wire n2217_o2_n;
  wire n2132_o2_p;
  wire n2132_o2_n;
  wire n2133_o2_p;
  wire n2133_o2_n;
  wire n2016_o2_p;
  wire n2016_o2_n;
  wire n2017_o2_p;
  wire n2017_o2_n;
  wire n1946_o2_p;
  wire n1946_o2_n;
  wire n1556_o2_p;
  wire n1556_o2_n;
  wire n1752_o2_p;
  wire n1752_o2_n;
  wire n1916_o2_p;
  wire n1916_o2_n;
  wire n2048_o2_p;
  wire n2048_o2_n;
  wire n2102_o2_p;
  wire n2102_o2_n;
  wire n1226_o2_p;
  wire n1226_o2_n;
  wire n1986_o2_p;
  wire n1986_o2_n;
  wire n1838_o2_p;
  wire n1838_o2_n;
  wire n1658_o2_p;
  wire n1658_o2_n;
  wire n829_inv_p;
  wire n829_inv_n;
  wire n1526_o2_p;
  wire n1526_o2_n;
  wire n1722_o2_p;
  wire n1722_o2_n;
  wire n1808_o2_p;
  wire n1808_o2_n;
  wire n1628_o2_p;
  wire n1628_o2_n;
  wire n844_inv_p;
  wire n844_inv_n;
  wire n847_inv_p;
  wire n847_inv_n;
  wire n1583_o2_p;
  wire n1583_o2_n;
  wire n1787_o2_p;
  wire n1787_o2_n;
  wire n1959_o2_p;
  wire n1959_o2_n;
  wire n2099_o2_p;
  wire n2099_o2_n;
  wire n2033_o2_p;
  wire n2033_o2_n;
  wire n1877_o2_p;
  wire n1877_o2_n;
  wire n1689_o2_p;
  wire n1689_o2_n;
  wire n1355_o2_p;
  wire n1355_o2_n;
  wire n1469_o2_p;
  wire n1469_o2_n;
  wire n1238_o2_p;
  wire n1238_o2_n;
  wire n1227_o2_p;
  wire n1227_o2_n;
  wire n1124_o2_p;
  wire n1124_o2_n;
  wire n704_o2_p;
  wire n704_o2_n;
  wire n484_o2_p;
  wire n484_o2_n;
  wire n1338_o2_p;
  wire n1338_o2_n;
  wire n1449_o2_p;
  wire n1449_o2_n;
  wire n1558_o2_p;
  wire n1558_o2_n;
  wire n1754_o2_p;
  wire n1754_o2_n;
  wire n1918_o2_p;
  wire n1918_o2_n;
  wire n2050_o2_p;
  wire n2050_o2_n;
  wire n2104_o2_p;
  wire n2104_o2_n;
  wire n1988_o2_p;
  wire n1988_o2_n;
  wire n1840_o2_p;
  wire n1840_o2_n;
  wire n1660_o2_p;
  wire n1660_o2_n;
  wire n708_o2_p;
  wire n708_o2_n;
  wire n768_o2_p;
  wire n768_o2_n;
  wire lo102_buf_o2_p;
  wire lo102_buf_o2_n;
  wire n1631_o2_p;
  wire n1631_o2_n;
  wire n1632_o2_p;
  wire n1632_o2_n;
  wire n1811_o2_p;
  wire n1811_o2_n;
  wire n1812_o2_p;
  wire n1812_o2_n;
  wire n1889_o2_p;
  wire n1889_o2_n;
  wire n1890_o2_p;
  wire n1890_o2_n;
  wire n1725_o2_p;
  wire n1725_o2_n;
  wire n1726_o2_p;
  wire n1726_o2_n;
  wire n917_o2_p;
  wire n917_o2_n;
  wire n918_o2_p;
  wire n918_o2_n;
  wire n1003_o2_p;
  wire n1003_o2_n;
  wire n1004_o2_p;
  wire n1004_o2_n;
  wire n1097_o2_p;
  wire n1097_o2_n;
  wire n1098_o2_p;
  wire n1098_o2_n;
  wire n1199_o2_p;
  wire n1199_o2_n;
  wire n1200_o2_p;
  wire n1200_o2_n;
  wire n1309_o2_p;
  wire n1309_o2_n;
  wire n1310_o2_p;
  wire n1310_o2_n;
  wire n1420_o2_p;
  wire n1420_o2_n;
  wire n1421_o2_p;
  wire n1421_o2_n;
  wire n1529_o2_p;
  wire n1529_o2_n;
  wire n1530_o2_p;
  wire n1530_o2_n;
  wire n839_o2_p;
  wire n839_o2_n;
  wire n840_o2_p;
  wire n840_o2_n;
  wire n577_o2_p;
  wire n577_o2_n;
  wire n623_o2_p;
  wire n623_o2_n;
  wire n677_o2_p;
  wire n677_o2_n;
  wire n739_o2_p;
  wire n739_o2_n;
  wire n809_o2_p;
  wire n809_o2_n;
  wire n887_o2_p;
  wire n887_o2_n;
  wire n973_o2_p;
  wire n973_o2_n;
  wire n1067_o2_p;
  wire n1067_o2_n;
  wire n1169_o2_p;
  wire n1169_o2_n;
  wire n1279_o2_p;
  wire n1279_o2_n;
  wire n1390_o2_p;
  wire n1390_o2_n;
  wire n1499_o2_p;
  wire n1499_o2_n;
  wire n539_o2_p;
  wire n539_o2_n;
  wire lo082_buf_o2_p;
  wire lo082_buf_o2_n;
  wire n555_o2_p;
  wire n555_o2_n;
  wire n601_o2_p;
  wire n601_o2_n;
  wire n655_o2_p;
  wire n655_o2_n;
  wire n717_o2_p;
  wire n717_o2_n;
  wire n787_o2_p;
  wire n787_o2_n;
  wire n865_o2_p;
  wire n865_o2_n;
  wire n951_o2_p;
  wire n951_o2_n;
  wire n1045_o2_p;
  wire n1045_o2_n;
  wire n1147_o2_p;
  wire n1147_o2_n;
  wire n1257_o2_p;
  wire n1257_o2_n;
  wire n1374_o2_p;
  wire n1374_o2_n;
  wire n1488_o2_p;
  wire n1488_o2_n;
  wire n1602_o2_p;
  wire n1602_o2_n;
  wire n517_o2_p;
  wire n517_o2_n;
  wire n1603_o2_p;
  wire n1603_o2_n;
  wire n509_o2_p;
  wire n509_o2_n;
  wire n510_o2_p;
  wire n510_o2_n;
  wire n579_o2_p;
  wire n579_o2_n;
  wire n625_o2_p;
  wire n625_o2_n;
  wire n679_o2_p;
  wire n679_o2_n;
  wire n741_o2_p;
  wire n741_o2_n;
  wire n811_o2_p;
  wire n811_o2_n;
  wire n889_o2_p;
  wire n889_o2_n;
  wire n975_o2_p;
  wire n975_o2_n;
  wire n1069_o2_p;
  wire n1069_o2_n;
  wire n1171_o2_p;
  wire n1171_o2_n;
  wire n1281_o2_p;
  wire n1281_o2_n;
  wire n1392_o2_p;
  wire n1392_o2_n;
  wire n1501_o2_p;
  wire n1501_o2_n;
  wire n541_o2_p;
  wire n541_o2_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire g1918_p;
  wire g1918_n;
  wire g1919_p;
  wire g1919_n;
  wire g1920_p;
  wire g1920_n;
  wire g1921_p;
  wire g1921_n;
  wire g1922_p;
  wire g1922_n;
  wire g1923_p;
  wire g1923_n;
  wire g1924_p;
  wire g1924_n;
  wire g1925_p;
  wire g1925_n;
  wire g1926_p;
  wire g1926_n;
  wire g1927_p;
  wire g1927_n;
  wire g1928_p;
  wire g1928_n;
  wire g1929_p;
  wire g1929_n;
  wire g1930_p;
  wire g1930_n;
  wire g1931_p;
  wire g1931_n;
  wire g1932_p;
  wire g1932_n;
  wire g1933_p;
  wire g1933_n;
  wire g1934_p;
  wire g1934_n;
  wire g1935_p;
  wire g1935_n;
  wire g1936_p;
  wire g1936_n;
  wire g1937_p;
  wire g1937_n;
  wire g1938_p;
  wire g1938_n;
  wire g1939_p;
  wire g1939_n;
  wire g1940_p;
  wire g1940_n;
  wire g1941_p;
  wire g1941_n;
  wire g1942_p;
  wire g1942_n;
  wire g1943_p;
  wire g1943_n;
  wire g1944_p;
  wire g1944_n;
  wire g1945_p;
  wire g1945_n;
  wire g1946_p;
  wire g1946_n;
  wire g1947_p;
  wire g1947_n;
  wire g1948_p;
  wire g1948_n;
  wire g1949_p;
  wire g1949_n;
  wire g1950_p;
  wire g1950_n;
  wire g1951_p;
  wire g1951_n;
  wire g1952_p;
  wire g1952_n;
  wire g1953_p;
  wire g1953_n;
  wire g1954_p;
  wire g1954_n;
  wire g1955_p;
  wire g1955_n;
  wire g1956_p;
  wire g1956_n;
  wire g1957_p;
  wire g1957_n;
  wire g1958_p;
  wire g1958_n;
  wire g1959_p;
  wire g1959_n;
  wire g1960_p;
  wire g1960_n;
  wire g1961_p;
  wire g1961_n;
  wire g1962_p;
  wire g1962_n;
  wire g1963_p;
  wire g1963_n;
  wire g1964_p;
  wire g1964_n;
  wire g1965_p;
  wire g1965_n;
  wire g1966_p;
  wire g1966_n;
  wire g1967_p;
  wire g1967_n;
  wire g1968_p;
  wire g1968_n;
  wire g1969_p;
  wire g1969_n;
  wire g1970_p;
  wire g1970_n;
  wire g1971_p;
  wire g1971_n;
  wire g1972_p;
  wire g1972_n;
  wire g1973_p;
  wire g1973_n;
  wire g1974_p;
  wire g1974_n;
  wire g1975_p;
  wire g1975_n;
  wire g1976_p;
  wire g1976_n;
  wire g1977_p;
  wire g1977_n;
  wire g1978_p;
  wire g1978_n;
  wire g1979_p;
  wire g1979_n;
  wire g1980_p;
  wire g1980_n;
  wire g1981_p;
  wire g1981_n;
  wire g1982_p;
  wire g1982_n;
  wire g1983_p;
  wire g1983_n;
  wire g1984_p;
  wire g1984_n;
  wire g1985_p;
  wire g1985_n;
  wire g1986_p;
  wire g1986_n;
  wire g1987_p;
  wire g1987_n;
  wire g1988_p;
  wire g1988_n;
  wire g1989_p;
  wire g1989_n;
  wire g1990_p;
  wire g1990_n;
  wire g1991_p;
  wire g1991_n;
  wire g1992_p;
  wire g1992_n;
  wire g1993_p;
  wire g1993_n;
  wire g1994_p;
  wire g1994_n;
  wire g1995_p;
  wire g1995_n;
  wire g1996_p;
  wire g1996_n;
  wire g1997_p;
  wire g1997_n;
  wire g1998_p;
  wire g1998_n;
  wire g1999_p;
  wire g1999_n;
  wire g2000_p;
  wire g2000_n;
  wire g2001_p;
  wire g2001_n;
  wire g2002_p;
  wire g2002_n;
  wire g2003_p;
  wire g2003_n;
  wire g2004_p;
  wire g2004_n;
  wire g2005_p;
  wire g2005_n;
  wire g2006_p;
  wire g2006_n;
  wire g2007_p;
  wire g2007_n;
  wire g2008_p;
  wire g2008_n;
  wire g2009_p;
  wire g2009_n;
  wire g2010_p;
  wire g2010_n;
  wire g2011_p;
  wire g2011_n;
  wire g2012_p;
  wire g2012_n;
  wire g2013_p;
  wire g2013_n;
  wire g2014_p;
  wire g2014_n;
  wire g2015_p;
  wire g2015_n;
  wire g2016_p;
  wire g2016_n;
  wire g2017_p;
  wire g2017_n;
  wire g2018_p;
  wire g2018_n;
  wire g2019_p;
  wire g2019_n;
  wire g2020_p;
  wire g2020_n;
  wire g2021_p;
  wire g2021_n;
  wire g2022_p;
  wire g2022_n;
  wire g2023_p;
  wire g2023_n;
  wire g2024_p;
  wire g2024_n;
  wire g2025_p;
  wire g2025_n;
  wire g2026_p;
  wire g2026_n;
  wire g2027_p;
  wire g2027_n;
  wire g2028_p;
  wire g2028_n;
  wire g2029_p;
  wire g2029_n;
  wire g2030_p;
  wire g2030_n;
  wire g2031_p;
  wire g2031_n;
  wire g2032_p;
  wire g2032_n;
  wire g2033_p;
  wire g2033_n;
  wire g2034_p;
  wire g2034_n;
  wire g2035_p;
  wire g2035_n;
  wire g2036_p;
  wire g2036_n;
  wire g2037_p;
  wire g2037_n;
  wire g2038_p;
  wire g2038_n;
  wire g2039_p;
  wire g2039_n;
  wire g2040_p;
  wire g2040_n;
  wire g2041_p;
  wire g2041_n;
  wire g2042_p;
  wire g2042_n;
  wire g2043_p;
  wire g2043_n;
  wire g2044_p;
  wire g2044_n;
  wire g2045_p;
  wire g2045_n;
  wire g2046_p;
  wire g2046_n;
  wire g2047_p;
  wire g2047_n;
  wire g2048_p;
  wire g2048_n;
  wire g2049_p;
  wire g2049_n;
  wire g2050_p;
  wire g2050_n;
  wire g2051_p;
  wire g2051_n;
  wire g2052_p;
  wire g2052_n;
  wire g2053_p;
  wire g2053_n;
  wire g2054_p;
  wire g2054_n;
  wire g2055_p;
  wire g2055_n;
  wire g2056_p;
  wire g2056_n;
  wire g2057_p;
  wire g2057_n;
  wire g2058_p;
  wire g2058_n;
  wire g2059_p;
  wire g2059_n;
  wire g2060_p;
  wire g2060_n;
  wire g2061_p;
  wire g2061_n;
  wire g2062_p;
  wire g2062_n;
  wire g2063_p;
  wire g2063_n;
  wire g2064_p;
  wire g2064_n;
  wire g2065_p;
  wire g2065_n;
  wire g2066_p;
  wire g2066_n;
  wire g2067_p;
  wire g2067_n;
  wire g2068_p;
  wire g2068_n;
  wire g2069_p;
  wire g2069_n;
  wire g2070_p;
  wire g2070_n;
  wire g2071_p;
  wire g2071_n;
  wire g2072_p;
  wire g2072_n;
  wire g2073_p;
  wire g2073_n;
  wire g2074_p;
  wire g2074_n;
  wire g2075_p;
  wire g2075_n;
  wire g2076_p;
  wire g2076_n;
  wire g2077_p;
  wire g2077_n;
  wire g2078_p;
  wire g2078_n;
  wire g2079_p;
  wire g2079_n;
  wire g2080_p;
  wire g2080_n;
  wire g2081_p;
  wire g2081_n;
  wire g2082_p;
  wire g2082_n;
  wire g2083_p;
  wire g2083_n;
  wire g2084_p;
  wire g2084_n;
  wire g2085_p;
  wire g2085_n;
  wire g2086_p;
  wire g2086_n;
  wire g2087_p;
  wire g2087_n;
  wire g2088_p;
  wire g2088_n;
  wire g2089_p;
  wire g2089_n;
  wire g2090_p;
  wire g2090_n;
  wire g2091_p;
  wire g2091_n;
  wire g2092_p;
  wire g2092_n;
  wire g2093_p;
  wire g2093_n;
  wire g2094_p;
  wire g2094_n;
  wire g2095_p;
  wire g2095_n;
  wire g2096_p;
  wire g2096_n;
  wire g2097_p;
  wire g2097_n;
  wire g2098_p;
  wire g2098_n;
  wire g2099_p;
  wire g2099_n;
  wire g2100_p;
  wire g2100_n;
  wire g2101_p;
  wire g2101_n;
  wire g2102_p;
  wire g2102_n;
  wire g2103_p;
  wire g2103_n;
  wire g2104_p;
  wire g2104_n;
  wire g2105_p;
  wire g2105_n;
  wire g2106_p;
  wire g2106_n;
  wire g2107_p;
  wire g2107_n;
  wire g2108_p;
  wire g2108_n;
  wire g2109_p;
  wire g2109_n;
  wire g2110_p;
  wire g2110_n;
  wire g2111_p;
  wire g2111_n;
  wire g2112_p;
  wire g2112_n;
  wire g2113_p;
  wire g2113_n;
  wire g2114_p;
  wire g2114_n;
  wire g2115_p;
  wire g2115_n;
  wire g2116_p;
  wire g2116_n;
  wire g2117_p;
  wire g2117_n;
  wire g2118_p;
  wire g2118_n;
  wire g2119_p;
  wire g2119_n;
  wire g2120_p;
  wire g2120_n;
  wire g2121_p;
  wire g2121_n;
  wire g2122_p;
  wire g2122_n;
  wire g2123_p;
  wire g2123_n;
  wire g2124_p;
  wire g2124_n;
  wire g2125_p;
  wire g2125_n;
  wire g2126_p;
  wire g2126_n;
  wire g2127_p;
  wire g2127_n;
  wire g2128_p;
  wire g2128_n;
  wire g2129_p;
  wire g2129_n;
  wire g2130_p;
  wire g2130_n;
  wire g2131_p;
  wire g2131_n;
  wire g2132_p;
  wire g2132_n;
  wire g2133_p;
  wire g2133_n;
  wire g2134_p;
  wire g2134_n;
  wire g2135_p;
  wire g2135_n;
  wire g2136_p;
  wire g2136_n;
  wire g2137_p;
  wire g2137_n;
  wire g2138_p;
  wire g2138_n;
  wire g2139_p;
  wire g2139_n;
  wire g2140_p;
  wire g2140_n;
  wire g2141_p;
  wire g2141_n;
  wire g2142_p;
  wire g2142_n;
  wire g2143_p;
  wire g2143_n;
  wire g2144_p;
  wire g2144_n;
  wire g2145_p;
  wire g2145_n;
  wire g2146_p;
  wire g2146_n;
  wire g2147_p;
  wire g2147_n;
  wire g2148_p;
  wire g2148_n;
  wire g2149_p;
  wire g2149_n;
  wire g2150_p;
  wire g2150_n;
  wire g2151_p;
  wire g2151_n;
  wire g2152_p;
  wire g2152_n;
  wire g2153_p;
  wire g2153_n;
  wire g2154_p;
  wire g2154_n;
  wire g2155_p;
  wire g2155_n;
  wire g2156_p;
  wire g2156_n;
  wire g2157_p;
  wire g2157_n;
  wire g2158_p;
  wire g2158_n;
  wire g2159_p;
  wire g2159_n;
  wire g2160_p;
  wire g2160_n;
  wire g2161_p;
  wire g2161_n;
  wire g2162_p;
  wire g2162_n;
  wire g2163_p;
  wire g2163_n;
  wire g2164_p;
  wire g2164_n;
  wire g2165_p;
  wire g2165_n;
  wire g2166_p;
  wire g2166_n;
  wire g2167_p;
  wire g2167_n;
  wire g2168_p;
  wire g2168_n;
  wire g2169_p;
  wire g2169_n;
  wire g2170_p;
  wire g2170_n;
  wire g2171_p;
  wire g2171_n;
  wire g2172_p;
  wire g2172_n;
  wire g2173_p;
  wire g2173_n;
  wire g2174_p;
  wire g2174_n;
  wire g2175_p;
  wire g2175_n;
  wire g2176_p;
  wire g2176_n;
  wire g2177_p;
  wire g2177_n;
  wire g2178_p;
  wire g2178_n;
  wire g2179_p;
  wire g2179_n;
  wire g2180_p;
  wire g2180_n;
  wire g2181_p;
  wire g2181_n;
  wire g2182_p;
  wire g2182_n;
  wire g2183_p;
  wire g2183_n;
  wire g2184_p;
  wire g2184_n;
  wire g2185_p;
  wire g2185_n;
  wire g2186_p;
  wire g2186_n;
  wire g2187_p;
  wire g2187_n;
  wire g2188_p;
  wire g2188_n;
  wire g2189_p;
  wire g2189_n;
  wire g2190_p;
  wire g2190_n;
  wire g2191_p;
  wire g2191_n;
  wire g2192_p;
  wire g2192_n;
  wire g2193_p;
  wire g2193_n;
  wire g2194_p;
  wire g2194_n;
  wire g2195_p;
  wire g2195_n;
  wire g2196_p;
  wire g2196_n;
  wire g2197_p;
  wire g2197_n;
  wire g2198_p;
  wire g2198_n;
  wire g2199_p;
  wire g2199_n;
  wire g2200_p;
  wire g2200_n;
  wire g2201_p;
  wire g2201_n;
  wire g2202_p;
  wire g2202_n;
  wire g2203_p;
  wire g2203_n;
  wire g2204_p;
  wire g2204_n;
  wire g2205_p;
  wire g2205_n;
  wire g2206_p;
  wire g2206_n;
  wire g2207_p;
  wire g2207_n;
  wire g2208_p;
  wire g2208_n;
  wire g2209_p;
  wire g2209_n;
  wire g2210_p;
  wire g2210_n;
  wire g2211_p;
  wire g2211_n;
  wire g2212_p;
  wire g2212_n;
  wire g2213_p;
  wire g2213_n;
  wire g2214_p;
  wire g2214_n;
  wire g2215_p;
  wire g2215_n;
  wire g2216_p;
  wire g2216_n;
  wire g2217_p;
  wire g2217_n;
  wire g2218_p;
  wire g2218_n;
  wire g2219_p;
  wire g2219_n;
  wire g2220_p;
  wire g2220_n;
  wire g2221_p;
  wire g2221_n;
  wire g2222_p;
  wire g2222_n;
  wire g2223_p;
  wire g2223_n;
  wire g2224_p;
  wire g2224_n;
  wire g2225_p;
  wire g2225_n;
  wire g2226_p;
  wire g2226_n;
  wire g2227_p;
  wire g2227_n;
  wire g2228_p;
  wire g2228_n;
  wire g2229_p;
  wire g2229_n;
  wire g2230_p;
  wire g2230_n;
  wire g2231_p;
  wire g2231_n;
  wire g2232_p;
  wire g2232_n;
  wire g2233_p;
  wire g2233_n;
  wire g2234_p;
  wire g2234_n;
  wire g2235_p;
  wire g2235_n;
  wire g2236_p;
  wire g2236_n;
  wire g2237_p;
  wire g2237_n;
  wire g2238_p;
  wire g2238_n;
  wire g2239_p;
  wire g2239_n;
  wire g2240_p;
  wire g2240_n;
  wire g2241_p;
  wire g2241_n;
  wire g2242_p;
  wire g2242_n;
  wire g2243_p;
  wire g2243_n;
  wire g2244_p;
  wire g2244_n;
  wire g2245_p;
  wire g2245_n;
  wire g2246_p;
  wire g2246_n;
  wire g2247_p;
  wire g2247_n;
  wire g2248_p;
  wire g2248_n;
  wire g2249_p;
  wire g2249_n;
  wire g2250_p;
  wire g2250_n;
  wire g2251_p;
  wire g2251_n;
  wire g2252_p;
  wire g2252_n;
  wire g2253_p;
  wire g2253_n;
  wire g2254_p;
  wire g2254_n;
  wire g2255_p;
  wire g2255_n;
  wire g2256_p;
  wire g2256_n;
  wire g2257_p;
  wire g2257_n;
  wire g2258_p;
  wire g2258_n;
  wire n1946_o2_p_spl_;
  wire n2016_o2_p_spl_;
  wire n2016_o2_n_spl_;
  wire g432_p_spl_;
  wire g433_n_spl_;
  wire g434_p_spl_;
  wire n2078_o2_n_spl_;
  wire n2078_o2_p_spl_;
  wire g438_n_spl_;
  wire g439_p_spl_;
  wire g438_p_spl_;
  wire g439_n_spl_;
  wire g440_n_spl_;
  wire g440_p_spl_;
  wire g437_p_spl_;
  wire g442_n_spl_;
  wire g443_p_spl_;
  wire n2863_lo_p_spl_;
  wire n2863_lo_p_spl_0;
  wire n2863_lo_p_spl_00;
  wire n2863_lo_p_spl_01;
  wire n2863_lo_p_spl_1;
  wire n2863_lo_p_spl_10;
  wire n2863_lo_n_spl_;
  wire n2863_lo_n_spl_0;
  wire n2863_lo_n_spl_00;
  wire n2863_lo_n_spl_01;
  wire n2863_lo_n_spl_1;
  wire n2863_lo_n_spl_10;
  wire n2132_o2_p_spl_;
  wire n2132_o2_n_spl_;
  wire g448_n_spl_;
  wire g449_p_spl_;
  wire g448_p_spl_;
  wire g449_n_spl_;
  wire g450_n_spl_;
  wire g450_p_spl_;
  wire g447_n_spl_;
  wire g452_p_spl_;
  wire g447_p_spl_;
  wire g452_n_spl_;
  wire g453_n_spl_;
  wire g453_p_spl_;
  wire g446_p_spl_;
  wire g455_n_spl_;
  wire g456_p_spl_;
  wire n2178_o2_n_spl_;
  wire n2178_o2_p_spl_;
  wire g462_n_spl_;
  wire g463_p_spl_;
  wire g462_p_spl_;
  wire g463_n_spl_;
  wire g464_n_spl_;
  wire g464_p_spl_;
  wire g461_n_spl_;
  wire g466_p_spl_;
  wire g461_p_spl_;
  wire g466_n_spl_;
  wire g467_n_spl_;
  wire g467_p_spl_;
  wire g460_n_spl_;
  wire g469_p_spl_;
  wire g460_p_spl_;
  wire g469_n_spl_;
  wire g470_n_spl_;
  wire g470_p_spl_;
  wire g459_p_spl_;
  wire g472_n_spl_;
  wire g473_p_spl_;
  wire n2635_lo_p_spl_;
  wire n2851_lo_p_spl_;
  wire n2851_lo_p_spl_0;
  wire n2851_lo_p_spl_1;
  wire n2635_lo_n_spl_;
  wire n2851_lo_n_spl_;
  wire n2851_lo_n_spl_0;
  wire n2851_lo_n_spl_1;
  wire n2216_o2_p_spl_;
  wire n2216_o2_n_spl_;
  wire g480_n_spl_;
  wire g481_p_spl_;
  wire g480_p_spl_;
  wire g481_n_spl_;
  wire g482_n_spl_;
  wire g482_p_spl_;
  wire g479_n_spl_;
  wire g484_p_spl_;
  wire g479_p_spl_;
  wire g484_n_spl_;
  wire g485_n_spl_;
  wire g485_p_spl_;
  wire g478_n_spl_;
  wire g487_p_spl_;
  wire g478_p_spl_;
  wire g487_n_spl_;
  wire g488_n_spl_;
  wire g488_p_spl_;
  wire g477_n_spl_;
  wire g490_p_spl_;
  wire g477_p_spl_;
  wire g490_n_spl_;
  wire g491_n_spl_;
  wire g491_p_spl_;
  wire g476_p_spl_;
  wire g493_n_spl_;
  wire g494_p_spl_;
  wire n2647_lo_p_spl_;
  wire n2647_lo_n_spl_;
  wire n2246_o2_n_spl_;
  wire n2246_o2_p_spl_;
  wire g502_n_spl_;
  wire g503_p_spl_;
  wire g502_p_spl_;
  wire g503_n_spl_;
  wire g504_n_spl_;
  wire g504_p_spl_;
  wire g501_n_spl_;
  wire g506_p_spl_;
  wire g501_p_spl_;
  wire g506_n_spl_;
  wire g507_n_spl_;
  wire g507_p_spl_;
  wire g500_n_spl_;
  wire g509_p_spl_;
  wire g500_p_spl_;
  wire g509_n_spl_;
  wire g510_n_spl_;
  wire g510_p_spl_;
  wire g499_n_spl_;
  wire g512_p_spl_;
  wire g499_p_spl_;
  wire g512_n_spl_;
  wire g513_n_spl_;
  wire g513_p_spl_;
  wire g498_n_spl_;
  wire g515_p_spl_;
  wire g498_p_spl_;
  wire g515_n_spl_;
  wire g516_n_spl_;
  wire g516_p_spl_;
  wire g497_p_spl_;
  wire g518_n_spl_;
  wire g519_p_spl_;
  wire n2659_lo_p_spl_;
  wire n2659_lo_n_spl_;
  wire n2671_lo_p_spl_;
  wire n2671_lo_p_spl_0;
  wire n2671_lo_n_spl_;
  wire n2671_lo_n_spl_0;
  wire g527_n_spl_;
  wire g528_n_spl_;
  wire g527_p_spl_;
  wire g528_p_spl_;
  wire g529_n_spl_;
  wire g529_p_spl_;
  wire g526_n_spl_;
  wire g531_p_spl_;
  wire g526_p_spl_;
  wire g531_n_spl_;
  wire g532_n_spl_;
  wire g532_p_spl_;
  wire g525_n_spl_;
  wire g534_p_spl_;
  wire g525_p_spl_;
  wire g534_n_spl_;
  wire g535_n_spl_;
  wire g535_p_spl_;
  wire g524_n_spl_;
  wire g537_p_spl_;
  wire g524_p_spl_;
  wire g537_n_spl_;
  wire g538_n_spl_;
  wire g538_p_spl_;
  wire g523_n_spl_;
  wire g540_p_spl_;
  wire g523_p_spl_;
  wire g540_n_spl_;
  wire g541_n_spl_;
  wire g541_p_spl_;
  wire g522_p_spl_;
  wire g543_n_spl_;
  wire g544_p_spl_;
  wire g550_n_spl_;
  wire g551_n_spl_;
  wire g550_p_spl_;
  wire g551_p_spl_;
  wire g552_n_spl_;
  wire g552_p_spl_;
  wire g549_n_spl_;
  wire g554_p_spl_;
  wire g549_p_spl_;
  wire g554_n_spl_;
  wire g555_n_spl_;
  wire g555_p_spl_;
  wire g548_n_spl_;
  wire g557_p_spl_;
  wire g548_p_spl_;
  wire g557_n_spl_;
  wire g558_n_spl_;
  wire g558_p_spl_;
  wire g547_p_spl_;
  wire g560_n_spl_;
  wire g561_p_spl_;
  wire g564_n_spl_;
  wire g565_n_spl_;
  wire g564_p_spl_;
  wire g565_p_spl_;
  wire g566_n_spl_;
  wire g570_n_spl_;
  wire n2848_lo_p_spl_;
  wire n2848_lo_p_spl_0;
  wire n2848_lo_p_spl_00;
  wire n2848_lo_p_spl_000;
  wire n2848_lo_p_spl_001;
  wire n2848_lo_p_spl_01;
  wire n2848_lo_p_spl_010;
  wire n2848_lo_p_spl_011;
  wire n2848_lo_p_spl_1;
  wire n2848_lo_p_spl_10;
  wire n2848_lo_p_spl_11;
  wire n4908_o2_p_spl_;
  wire n2848_lo_n_spl_;
  wire n2848_lo_n_spl_0;
  wire n2848_lo_n_spl_00;
  wire n2848_lo_n_spl_000;
  wire n2848_lo_n_spl_001;
  wire n2848_lo_n_spl_01;
  wire n2848_lo_n_spl_010;
  wire n2848_lo_n_spl_011;
  wire n2848_lo_n_spl_1;
  wire n2848_lo_n_spl_10;
  wire n2848_lo_n_spl_11;
  wire n4908_o2_n_spl_;
  wire n1124_o2_p_spl_;
  wire g575_n_spl_;
  wire g576_p_spl_;
  wire g575_p_spl_;
  wire g576_n_spl_;
  wire g577_n_spl_;
  wire g577_p_spl_;
  wire g579_p_spl_;
  wire g574_p_spl_;
  wire n2860_lo_n_spl_;
  wire n2860_lo_n_spl_0;
  wire n2860_lo_n_spl_00;
  wire n2860_lo_n_spl_000;
  wire n2860_lo_n_spl_01;
  wire n2860_lo_n_spl_1;
  wire n2860_lo_n_spl_10;
  wire n2860_lo_n_spl_11;
  wire g580_p_spl_;
  wire n4867_o2_p_spl_;
  wire n4867_o2_n_spl_;
  wire n1238_o2_n_spl_;
  wire n1338_o2_n_spl_;
  wire n1238_o2_p_spl_;
  wire n1338_o2_p_spl_;
  wire g584_n_spl_;
  wire g584_p_spl_;
  wire g583_n_spl_;
  wire g586_p_spl_;
  wire g583_p_spl_;
  wire g586_n_spl_;
  wire g587_n_spl_;
  wire g587_p_spl_;
  wire g582_n_spl_;
  wire g589_p_spl_;
  wire g581_n_spl_;
  wire g592_p_spl_;
  wire g593_p_spl_;
  wire n2860_lo_p_spl_;
  wire n2860_lo_p_spl_0;
  wire n2860_lo_p_spl_00;
  wire n2860_lo_p_spl_01;
  wire n2860_lo_p_spl_1;
  wire n2860_lo_p_spl_10;
  wire n2860_lo_p_spl_11;
  wire n4836_o2_p_spl_;
  wire n4836_o2_n_spl_;
  wire n1355_o2_n_spl_;
  wire n1449_o2_n_spl_;
  wire n1355_o2_p_spl_;
  wire n1449_o2_p_spl_;
  wire g598_n_spl_;
  wire g598_p_spl_;
  wire g597_n_spl_;
  wire g600_p_spl_;
  wire g597_p_spl_;
  wire g600_n_spl_;
  wire g601_n_spl_;
  wire g601_p_spl_;
  wire g596_n_spl_;
  wire g603_p_spl_;
  wire g596_p_spl_;
  wire g603_n_spl_;
  wire g604_n_spl_;
  wire g604_p_spl_;
  wire g595_n_spl_;
  wire g606_p_spl_;
  wire g607_n_spl_;
  wire g594_n_spl_;
  wire g609_p_spl_;
  wire n4837_o2_p_spl_;
  wire n4837_o2_n_spl_;
  wire n1469_o2_n_spl_;
  wire n1558_o2_n_spl_;
  wire n1469_o2_p_spl_;
  wire n1558_o2_p_spl_;
  wire g615_n_spl_;
  wire g615_p_spl_;
  wire g614_n_spl_;
  wire g617_p_spl_;
  wire g614_p_spl_;
  wire g617_n_spl_;
  wire g618_n_spl_;
  wire g618_p_spl_;
  wire g613_n_spl_;
  wire g620_p_spl_;
  wire g613_p_spl_;
  wire g620_n_spl_;
  wire g621_n_spl_;
  wire g621_p_spl_;
  wire g612_n_spl_;
  wire g623_p_spl_;
  wire g612_p_spl_;
  wire g623_n_spl_;
  wire g624_n_spl_;
  wire g624_p_spl_;
  wire g611_n_spl_;
  wire g626_p_spl_;
  wire n6148_o2_p_spl_;
  wire n6148_o2_p_spl_0;
  wire n6148_o2_p_spl_00;
  wire n6148_o2_p_spl_1;
  wire lo102_buf_o2_p_spl_;
  wire lo102_buf_o2_p_spl_0;
  wire lo102_buf_o2_p_spl_00;
  wire lo102_buf_o2_p_spl_000;
  wire lo102_buf_o2_p_spl_001;
  wire lo102_buf_o2_p_spl_01;
  wire lo102_buf_o2_p_spl_010;
  wire lo102_buf_o2_p_spl_011;
  wire lo102_buf_o2_p_spl_1;
  wire lo102_buf_o2_p_spl_10;
  wire lo102_buf_o2_p_spl_100;
  wire lo102_buf_o2_p_spl_101;
  wire lo102_buf_o2_p_spl_11;
  wire lo102_buf_o2_p_spl_110;
  wire lo102_buf_o2_p_spl_111;
  wire n6148_o2_n_spl_;
  wire n6148_o2_n_spl_0;
  wire n6148_o2_n_spl_00;
  wire n6148_o2_n_spl_1;
  wire lo102_buf_o2_n_spl_;
  wire lo102_buf_o2_n_spl_0;
  wire lo102_buf_o2_n_spl_00;
  wire lo102_buf_o2_n_spl_000;
  wire lo102_buf_o2_n_spl_001;
  wire lo102_buf_o2_n_spl_01;
  wire lo102_buf_o2_n_spl_010;
  wire lo102_buf_o2_n_spl_011;
  wire lo102_buf_o2_n_spl_1;
  wire lo102_buf_o2_n_spl_10;
  wire lo102_buf_o2_n_spl_100;
  wire lo102_buf_o2_n_spl_101;
  wire lo102_buf_o2_n_spl_11;
  wire lo102_buf_o2_n_spl_110;
  wire lo102_buf_o2_n_spl_111;
  wire g610_n_spl_;
  wire g629_p_spl_;
  wire n708_o2_n_spl_;
  wire n768_o2_n_spl_;
  wire n708_o2_p_spl_;
  wire n768_o2_p_spl_;
  wire g632_n_spl_;
  wire g632_p_spl_;
  wire g634_p_spl_;
  wire g630_p_spl_;
  wire g631_p_spl_;
  wire n4838_o2_p_spl_;
  wire n4838_o2_n_spl_;
  wire n1583_o2_n_spl_;
  wire n1660_o2_p_spl_;
  wire n1583_o2_p_spl_;
  wire n1660_o2_n_spl_;
  wire g642_n_spl_;
  wire g642_p_spl_;
  wire g641_n_spl_;
  wire g644_p_spl_;
  wire g641_p_spl_;
  wire g644_n_spl_;
  wire g645_n_spl_;
  wire g645_p_spl_;
  wire g640_n_spl_;
  wire g647_p_spl_;
  wire g640_p_spl_;
  wire g647_n_spl_;
  wire g648_n_spl_;
  wire g648_p_spl_;
  wire g639_n_spl_;
  wire g650_p_spl_;
  wire g639_p_spl_;
  wire g650_n_spl_;
  wire g651_n_spl_;
  wire g651_p_spl_;
  wire g638_n_spl_;
  wire g653_p_spl_;
  wire g638_p_spl_;
  wire g653_n_spl_;
  wire g654_n_spl_;
  wire g654_p_spl_;
  wire g637_n_spl_;
  wire g656_p_spl_;
  wire n2797_lo_p_spl_;
  wire n2797_lo_p_spl_0;
  wire n2797_lo_p_spl_00;
  wire n2797_lo_p_spl_000;
  wire n2797_lo_p_spl_001;
  wire n2797_lo_p_spl_01;
  wire n2797_lo_p_spl_010;
  wire n2797_lo_p_spl_011;
  wire n2797_lo_p_spl_1;
  wire n2797_lo_p_spl_10;
  wire n2797_lo_p_spl_100;
  wire n2797_lo_p_spl_101;
  wire n2797_lo_p_spl_11;
  wire n2797_lo_p_spl_110;
  wire n2797_lo_p_spl_111;
  wire n2797_lo_n_spl_;
  wire n2797_lo_n_spl_0;
  wire n2797_lo_n_spl_00;
  wire n2797_lo_n_spl_000;
  wire n2797_lo_n_spl_001;
  wire n2797_lo_n_spl_01;
  wire n2797_lo_n_spl_010;
  wire n2797_lo_n_spl_011;
  wire n2797_lo_n_spl_1;
  wire n2797_lo_n_spl_10;
  wire n2797_lo_n_spl_100;
  wire n2797_lo_n_spl_101;
  wire n2797_lo_n_spl_11;
  wire g636_n_spl_;
  wire g659_p_spl_;
  wire g635_p_spl_;
  wire n6053_o2_p_spl_;
  wire n6053_o2_p_spl_0;
  wire n6053_o2_p_spl_00;
  wire n6053_o2_p_spl_1;
  wire n6053_o2_n_spl_;
  wire n6053_o2_n_spl_0;
  wire n6053_o2_n_spl_00;
  wire n6053_o2_n_spl_1;
  wire n839_o2_p_spl_;
  wire n839_o2_n_spl_;
  wire g663_n_spl_;
  wire g664_p_spl_;
  wire g663_p_spl_;
  wire g664_n_spl_;
  wire g665_n_spl_;
  wire g665_p_spl_;
  wire g662_n_spl_;
  wire g667_p_spl_;
  wire g662_p_spl_;
  wire g667_n_spl_;
  wire g668_n_spl_;
  wire g668_p_spl_;
  wire g670_p_spl_;
  wire g660_p_spl_;
  wire lo002_buf_o2_p_spl_;
  wire lo002_buf_o2_p_spl_0;
  wire lo002_buf_o2_p_spl_00;
  wire lo002_buf_o2_p_spl_1;
  wire lo082_buf_o2_p_spl_;
  wire lo082_buf_o2_p_spl_0;
  wire lo002_buf_o2_n_spl_;
  wire lo002_buf_o2_n_spl_0;
  wire lo002_buf_o2_n_spl_00;
  wire lo002_buf_o2_n_spl_1;
  wire lo082_buf_o2_n_spl_;
  wire lo082_buf_o2_n_spl_0;
  wire n509_o2_p_spl_;
  wire n509_o2_n_spl_;
  wire g661_p_spl_;
  wire n4839_o2_p_spl_;
  wire n4839_o2_n_spl_;
  wire n4840_o2_p_spl_;
  wire n4840_o2_p_spl_0;
  wire lo118_buf_o2_p_spl_;
  wire lo118_buf_o2_p_spl_0;
  wire lo118_buf_o2_p_spl_00;
  wire lo118_buf_o2_p_spl_000;
  wire lo118_buf_o2_p_spl_01;
  wire lo118_buf_o2_p_spl_1;
  wire lo118_buf_o2_p_spl_10;
  wire lo118_buf_o2_p_spl_11;
  wire n4840_o2_n_spl_;
  wire n4840_o2_n_spl_0;
  wire lo118_buf_o2_n_spl_;
  wire lo118_buf_o2_n_spl_0;
  wire lo118_buf_o2_n_spl_00;
  wire lo118_buf_o2_n_spl_000;
  wire lo118_buf_o2_n_spl_01;
  wire lo118_buf_o2_n_spl_1;
  wire lo118_buf_o2_n_spl_10;
  wire lo118_buf_o2_n_spl_11;
  wire n1689_o2_n_spl_;
  wire n1754_o2_n_spl_;
  wire n1689_o2_p_spl_;
  wire n1754_o2_p_spl_;
  wire g681_n_spl_;
  wire g681_p_spl_;
  wire g680_n_spl_;
  wire g683_p_spl_;
  wire g680_p_spl_;
  wire g683_n_spl_;
  wire g684_n_spl_;
  wire g684_p_spl_;
  wire g679_n_spl_;
  wire g686_p_spl_;
  wire g679_p_spl_;
  wire g686_n_spl_;
  wire g687_n_spl_;
  wire g687_p_spl_;
  wire g678_n_spl_;
  wire g689_p_spl_;
  wire g678_p_spl_;
  wire g689_n_spl_;
  wire g690_n_spl_;
  wire g690_p_spl_;
  wire g677_n_spl_;
  wire g692_p_spl_;
  wire g677_p_spl_;
  wire g692_n_spl_;
  wire g693_n_spl_;
  wire g693_p_spl_;
  wire g676_n_spl_;
  wire g695_p_spl_;
  wire g676_p_spl_;
  wire g695_n_spl_;
  wire g696_n_spl_;
  wire g696_p_spl_;
  wire g675_n_spl_;
  wire g698_p_spl_;
  wire g673_p_spl_;
  wire g672_p_spl_;
  wire n2809_lo_p_spl_;
  wire n2809_lo_p_spl_0;
  wire n2809_lo_p_spl_00;
  wire n2809_lo_p_spl_000;
  wire n2809_lo_p_spl_001;
  wire n2809_lo_p_spl_01;
  wire n2809_lo_p_spl_010;
  wire n2809_lo_p_spl_011;
  wire n2809_lo_p_spl_1;
  wire n2809_lo_p_spl_10;
  wire n2809_lo_p_spl_100;
  wire n2809_lo_p_spl_11;
  wire n2809_lo_n_spl_;
  wire n2809_lo_n_spl_0;
  wire n2809_lo_n_spl_00;
  wire n2809_lo_n_spl_000;
  wire n2809_lo_n_spl_001;
  wire n2809_lo_n_spl_01;
  wire n2809_lo_n_spl_010;
  wire n2809_lo_n_spl_1;
  wire n2809_lo_n_spl_10;
  wire n2809_lo_n_spl_11;
  wire n2734_lo_p_spl_;
  wire n2734_lo_p_spl_0;
  wire n2734_lo_p_spl_00;
  wire n2734_lo_p_spl_000;
  wire n2734_lo_p_spl_001;
  wire n2734_lo_p_spl_01;
  wire n2734_lo_p_spl_010;
  wire n2734_lo_p_spl_011;
  wire n2734_lo_p_spl_1;
  wire n2734_lo_p_spl_10;
  wire n2734_lo_p_spl_100;
  wire n2734_lo_p_spl_101;
  wire n2734_lo_p_spl_11;
  wire n2734_lo_p_spl_110;
  wire n2734_lo_p_spl_111;
  wire n2734_lo_n_spl_;
  wire n2734_lo_n_spl_0;
  wire n2734_lo_n_spl_00;
  wire n2734_lo_n_spl_000;
  wire n2734_lo_n_spl_001;
  wire n2734_lo_n_spl_01;
  wire n2734_lo_n_spl_010;
  wire n2734_lo_n_spl_011;
  wire n2734_lo_n_spl_1;
  wire n2734_lo_n_spl_10;
  wire n2734_lo_n_spl_100;
  wire n2734_lo_n_spl_101;
  wire n2734_lo_n_spl_11;
  wire n2734_lo_n_spl_110;
  wire n2734_lo_n_spl_111;
  wire n2099_o2_n_spl_;
  wire n2104_o2_p_spl_;
  wire n2099_o2_p_spl_;
  wire n2104_o2_n_spl_;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire g705_n_spl_;
  wire g708_p_spl_;
  wire g705_p_spl_;
  wire g708_n_spl_;
  wire n4847_o2_p_spl_;
  wire n4847_o2_p_spl_0;
  wire n4847_o2_p_spl_1;
  wire lo110_buf_o2_p_spl_;
  wire lo110_buf_o2_p_spl_0;
  wire lo110_buf_o2_p_spl_1;
  wire n4847_o2_n_spl_;
  wire n4847_o2_n_spl_0;
  wire lo110_buf_o2_n_spl_;
  wire lo110_buf_o2_n_spl_0;
  wire lo110_buf_o2_n_spl_1;
  wire g709_n_spl_;
  wire g709_p_spl_;
  wire g710_n_spl_;
  wire g712_p_spl_;
  wire g710_p_spl_;
  wire g712_n_spl_;
  wire g713_n_spl_;
  wire g713_p_spl_;
  wire n4848_o2_p_spl_;
  wire n4848_o2_p_spl_0;
  wire n4848_o2_n_spl_;
  wire n4848_o2_n_spl_0;
  wire n4849_o2_p_spl_;
  wire n4849_o2_p_spl_0;
  wire n4849_o2_p_spl_1;
  wire n4849_o2_n_spl_;
  wire n4849_o2_n_spl_0;
  wire g716_n_spl_;
  wire g717_n_spl_;
  wire g716_p_spl_;
  wire g717_p_spl_;
  wire g718_n_spl_;
  wire g718_p_spl_;
  wire g715_n_spl_;
  wire g720_p_spl_;
  wire g715_p_spl_;
  wire g720_n_spl_;
  wire g721_n_spl_;
  wire g721_p_spl_;
  wire g714_n_spl_;
  wire g723_p_spl_;
  wire g714_p_spl_;
  wire g723_n_spl_;
  wire lo114_buf_o2_p_spl_;
  wire lo114_buf_o2_p_spl_0;
  wire lo114_buf_o2_p_spl_00;
  wire lo114_buf_o2_p_spl_01;
  wire lo114_buf_o2_p_spl_1;
  wire lo114_buf_o2_p_spl_10;
  wire lo114_buf_o2_n_spl_;
  wire lo114_buf_o2_n_spl_0;
  wire lo114_buf_o2_n_spl_00;
  wire lo114_buf_o2_n_spl_01;
  wire lo114_buf_o2_n_spl_1;
  wire lo114_buf_o2_n_spl_10;
  wire g724_n_spl_;
  wire g724_p_spl_;
  wire g725_n_spl_;
  wire g727_p_spl_;
  wire g725_p_spl_;
  wire g727_n_spl_;
  wire g728_n_spl_;
  wire g728_p_spl_;
  wire g731_n_spl_;
  wire g732_n_spl_;
  wire g731_p_spl_;
  wire g732_p_spl_;
  wire g733_n_spl_;
  wire g733_p_spl_;
  wire g730_n_spl_;
  wire g735_p_spl_;
  wire g730_p_spl_;
  wire g735_n_spl_;
  wire g736_n_spl_;
  wire g736_p_spl_;
  wire g729_n_spl_;
  wire g738_p_spl_;
  wire g729_p_spl_;
  wire g738_n_spl_;
  wire n1959_o2_n_spl_;
  wire n1988_o2_p_spl_;
  wire n1959_o2_p_spl_;
  wire n1988_o2_n_spl_;
  wire g741_n_spl_;
  wire g741_p_spl_;
  wire g740_n_spl_;
  wire g743_p_spl_;
  wire g740_p_spl_;
  wire g743_n_spl_;
  wire n4844_o2_p_spl_;
  wire n4844_o2_p_spl_0;
  wire n4844_o2_p_spl_1;
  wire n4844_o2_n_spl_;
  wire n4844_o2_n_spl_0;
  wire g744_n_spl_;
  wire g744_p_spl_;
  wire g745_n_spl_;
  wire g747_p_spl_;
  wire g745_p_spl_;
  wire g747_n_spl_;
  wire g748_n_spl_;
  wire g748_p_spl_;
  wire n4845_o2_p_spl_;
  wire n4845_o2_p_spl_0;
  wire n4845_o2_n_spl_;
  wire n4845_o2_n_spl_0;
  wire n4846_o2_p_spl_;
  wire n4846_o2_p_spl_0;
  wire n4846_o2_p_spl_1;
  wire n4846_o2_n_spl_;
  wire n4846_o2_n_spl_0;
  wire n2033_o2_n_spl_;
  wire n2050_o2_n_spl_;
  wire n2033_o2_p_spl_;
  wire n2050_o2_p_spl_;
  wire g753_n_spl_;
  wire g753_p_spl_;
  wire g752_n_spl_;
  wire g755_p_spl_;
  wire g752_p_spl_;
  wire g755_n_spl_;
  wire g756_n_spl_;
  wire g756_p_spl_;
  wire g751_n_spl_;
  wire g758_p_spl_;
  wire g751_p_spl_;
  wire g758_n_spl_;
  wire g759_n_spl_;
  wire g759_p_spl_;
  wire g750_n_spl_;
  wire g761_p_spl_;
  wire g750_p_spl_;
  wire g761_n_spl_;
  wire g762_n_spl_;
  wire g762_p_spl_;
  wire g749_n_spl_;
  wire g764_p_spl_;
  wire g749_p_spl_;
  wire g764_n_spl_;
  wire g765_n_spl_;
  wire g765_p_spl_;
  wire g766_n_spl_;
  wire g768_p_spl_;
  wire g766_p_spl_;
  wire g768_n_spl_;
  wire g769_n_spl_;
  wire g769_p_spl_;
  wire g774_n_spl_;
  wire g776_p_spl_;
  wire g774_p_spl_;
  wire g776_n_spl_;
  wire g777_n_spl_;
  wire g777_p_spl_;
  wire g773_n_spl_;
  wire g779_p_spl_;
  wire g773_p_spl_;
  wire g779_n_spl_;
  wire g780_n_spl_;
  wire g780_p_spl_;
  wire g772_n_spl_;
  wire g782_p_spl_;
  wire g772_p_spl_;
  wire g782_n_spl_;
  wire g783_n_spl_;
  wire g783_p_spl_;
  wire g771_n_spl_;
  wire g785_p_spl_;
  wire g771_p_spl_;
  wire g785_n_spl_;
  wire g786_n_spl_;
  wire g786_p_spl_;
  wire g770_n_spl_;
  wire g788_p_spl_;
  wire g770_p_spl_;
  wire g788_n_spl_;
  wire n1787_o2_n_spl_;
  wire n1840_o2_p_spl_;
  wire n1787_o2_p_spl_;
  wire n1840_o2_n_spl_;
  wire g791_n_spl_;
  wire g791_p_spl_;
  wire g790_n_spl_;
  wire g793_p_spl_;
  wire g790_p_spl_;
  wire g793_n_spl_;
  wire n4841_o2_p_spl_;
  wire n4841_o2_p_spl_0;
  wire n4841_o2_n_spl_;
  wire n4841_o2_n_spl_0;
  wire g794_n_spl_;
  wire g794_p_spl_;
  wire g795_n_spl_;
  wire g797_p_spl_;
  wire g795_p_spl_;
  wire g797_n_spl_;
  wire g798_n_spl_;
  wire g798_p_spl_;
  wire n4842_o2_p_spl_;
  wire n4842_o2_n_spl_;
  wire n4842_o2_n_spl_0;
  wire n4843_o2_p_spl_;
  wire n4843_o2_p_spl_0;
  wire n4843_o2_p_spl_1;
  wire n4843_o2_n_spl_;
  wire n4843_o2_n_spl_0;
  wire n1877_o2_n_spl_;
  wire n1918_o2_n_spl_;
  wire n1877_o2_p_spl_;
  wire n1918_o2_p_spl_;
  wire g803_n_spl_;
  wire g803_p_spl_;
  wire g802_n_spl_;
  wire g805_p_spl_;
  wire g802_p_spl_;
  wire g805_n_spl_;
  wire g806_n_spl_;
  wire g806_p_spl_;
  wire g801_n_spl_;
  wire g808_p_spl_;
  wire g801_p_spl_;
  wire g808_n_spl_;
  wire g809_n_spl_;
  wire g809_p_spl_;
  wire g800_n_spl_;
  wire g811_p_spl_;
  wire g800_p_spl_;
  wire g811_n_spl_;
  wire g812_n_spl_;
  wire g812_p_spl_;
  wire g799_n_spl_;
  wire g814_p_spl_;
  wire g799_p_spl_;
  wire g814_n_spl_;
  wire g815_n_spl_;
  wire g815_p_spl_;
  wire g816_n_spl_;
  wire g818_p_spl_;
  wire g816_p_spl_;
  wire g818_n_spl_;
  wire g819_n_spl_;
  wire g819_p_spl_;
  wire g824_n_spl_;
  wire g826_p_spl_;
  wire g824_p_spl_;
  wire g826_n_spl_;
  wire g827_n_spl_;
  wire g827_p_spl_;
  wire g823_n_spl_;
  wire g829_p_spl_;
  wire g823_p_spl_;
  wire g829_n_spl_;
  wire g830_n_spl_;
  wire g830_p_spl_;
  wire g822_n_spl_;
  wire g832_p_spl_;
  wire g822_p_spl_;
  wire g832_n_spl_;
  wire g833_n_spl_;
  wire g833_p_spl_;
  wire g821_n_spl_;
  wire g835_p_spl_;
  wire g821_p_spl_;
  wire g835_n_spl_;
  wire g836_n_spl_;
  wire g836_p_spl_;
  wire g820_n_spl_;
  wire g838_p_spl_;
  wire g820_p_spl_;
  wire g838_n_spl_;
  wire g674_n_spl_;
  wire g701_p_spl_;
  wire g671_p_spl_;
  wire n6024_o2_p_spl_;
  wire n6024_o2_p_spl_0;
  wire n6024_o2_p_spl_00;
  wire n6024_o2_p_spl_01;
  wire n6024_o2_p_spl_1;
  wire n6024_o2_n_spl_;
  wire n6024_o2_n_spl_0;
  wire n6024_o2_n_spl_00;
  wire n6024_o2_n_spl_1;
  wire n917_o2_p_spl_;
  wire n917_o2_n_spl_;
  wire g844_n_spl_;
  wire g845_p_spl_;
  wire g844_p_spl_;
  wire g845_n_spl_;
  wire g846_n_spl_;
  wire g846_p_spl_;
  wire g843_n_spl_;
  wire g848_p_spl_;
  wire g843_p_spl_;
  wire g848_n_spl_;
  wire g849_n_spl_;
  wire g849_p_spl_;
  wire g842_n_spl_;
  wire g851_p_spl_;
  wire g842_p_spl_;
  wire g851_n_spl_;
  wire g852_n_spl_;
  wire g852_p_spl_;
  wire g841_n_spl_;
  wire g854_p_spl_;
  wire g841_p_spl_;
  wire g854_n_spl_;
  wire g855_n_spl_;
  wire g855_p_spl_;
  wire g702_p_spl_;
  wire n517_o2_n_spl_;
  wire n541_o2_p_spl_;
  wire n517_o2_p_spl_;
  wire n541_o2_n_spl_;
  wire g859_n_spl_;
  wire g859_p_spl_;
  wire g858_n_spl_;
  wire g861_p_spl_;
  wire g858_p_spl_;
  wire g861_n_spl_;
  wire g862_n_spl_;
  wire g862_p_spl_;
  wire g857_p_spl_;
  wire g703_p_spl_;
  wire g864_p_spl_;
  wire g704_p_spl_;
  wire g840_p_spl_;
  wire g872_n_spl_;
  wire g874_p_spl_;
  wire g872_p_spl_;
  wire g874_n_spl_;
  wire g875_n_spl_;
  wire g875_p_spl_;
  wire g871_n_spl_;
  wire g877_p_spl_;
  wire g871_p_spl_;
  wire g877_n_spl_;
  wire g878_n_spl_;
  wire g878_p_spl_;
  wire g870_n_spl_;
  wire g880_p_spl_;
  wire g870_p_spl_;
  wire g880_n_spl_;
  wire g881_n_spl_;
  wire g881_p_spl_;
  wire g869_n_spl_;
  wire g883_p_spl_;
  wire g869_p_spl_;
  wire g883_n_spl_;
  wire g884_n_spl_;
  wire g884_p_spl_;
  wire g868_n_spl_;
  wire g886_p_spl_;
  wire n2746_lo_p_spl_;
  wire n2746_lo_p_spl_0;
  wire n2746_lo_p_spl_00;
  wire n2746_lo_p_spl_000;
  wire n2746_lo_p_spl_001;
  wire n2746_lo_p_spl_01;
  wire n2746_lo_p_spl_010;
  wire n2746_lo_p_spl_011;
  wire n2746_lo_p_spl_1;
  wire n2746_lo_p_spl_10;
  wire n2746_lo_p_spl_100;
  wire n2746_lo_p_spl_101;
  wire n2746_lo_p_spl_11;
  wire n2746_lo_p_spl_110;
  wire n2746_lo_n_spl_;
  wire n2746_lo_n_spl_0;
  wire n2746_lo_n_spl_00;
  wire n2746_lo_n_spl_000;
  wire n2746_lo_n_spl_001;
  wire n2746_lo_n_spl_01;
  wire n2746_lo_n_spl_010;
  wire n2746_lo_n_spl_011;
  wire n2746_lo_n_spl_1;
  wire n2746_lo_n_spl_10;
  wire n2746_lo_n_spl_100;
  wire n2746_lo_n_spl_101;
  wire n2746_lo_n_spl_11;
  wire n2746_lo_n_spl_110;
  wire n2746_lo_n_spl_111;
  wire g866_p_spl_;
  wire lo006_buf_o2_p_spl_;
  wire lo006_buf_o2_p_spl_0;
  wire lo006_buf_o2_p_spl_00;
  wire lo006_buf_o2_p_spl_1;
  wire lo006_buf_o2_n_spl_;
  wire lo006_buf_o2_n_spl_0;
  wire lo006_buf_o2_n_spl_1;
  wire n555_o2_n_spl_;
  wire n579_o2_p_spl_;
  wire n555_o2_p_spl_;
  wire n579_o2_n_spl_;
  wire g894_n_spl_;
  wire g894_p_spl_;
  wire g893_n_spl_;
  wire g896_p_spl_;
  wire g893_p_spl_;
  wire g896_n_spl_;
  wire g897_n_spl_;
  wire g897_p_spl_;
  wire g892_n_spl_;
  wire g899_p_spl_;
  wire g892_p_spl_;
  wire g899_n_spl_;
  wire g900_n_spl_;
  wire g900_p_spl_;
  wire g891_n_spl_;
  wire g902_p_spl_;
  wire g891_p_spl_;
  wire g902_n_spl_;
  wire g903_n_spl_;
  wire g903_p_spl_;
  wire g905_p_spl_;
  wire g890_p_spl_;
  wire n2821_lo_p_spl_;
  wire n2821_lo_p_spl_0;
  wire n2821_lo_p_spl_00;
  wire n2821_lo_p_spl_000;
  wire n2821_lo_p_spl_001;
  wire n2821_lo_p_spl_01;
  wire n2821_lo_p_spl_1;
  wire n2821_lo_p_spl_10;
  wire n2821_lo_p_spl_11;
  wire n2821_lo_n_spl_;
  wire n2821_lo_n_spl_0;
  wire n2821_lo_n_spl_00;
  wire n2821_lo_n_spl_01;
  wire n2821_lo_n_spl_1;
  wire n2821_lo_n_spl_10;
  wire n2821_lo_n_spl_11;
  wire g839_n_spl_;
  wire g789_n_spl_;
  wire g739_n_spl_;
  wire g925_n_spl_;
  wire g927_p_spl_;
  wire g925_p_spl_;
  wire g927_n_spl_;
  wire g928_p_spl_;
  wire g924_n_spl_;
  wire g930_p_spl_;
  wire g924_p_spl_;
  wire g930_n_spl_;
  wire g931_p_spl_;
  wire g937_n_spl_;
  wire g939_p_spl_;
  wire g937_p_spl_;
  wire g939_n_spl_;
  wire g940_p_spl_;
  wire g936_n_spl_;
  wire g942_p_spl_;
  wire g936_p_spl_;
  wire g942_n_spl_;
  wire g943_p_spl_;
  wire g949_n_spl_;
  wire g951_p_spl_;
  wire g949_p_spl_;
  wire g951_n_spl_;
  wire g952_p_spl_;
  wire g948_n_spl_;
  wire g954_p_spl_;
  wire g948_p_spl_;
  wire g954_n_spl_;
  wire g955_p_spl_;
  wire g867_n_spl_;
  wire g889_p_spl_;
  wire g865_p_spl_;
  wire n6025_o2_p_spl_;
  wire n6025_o2_p_spl_0;
  wire n6025_o2_p_spl_00;
  wire n6025_o2_p_spl_01;
  wire n6025_o2_p_spl_1;
  wire n6025_o2_n_spl_;
  wire n6025_o2_n_spl_0;
  wire n6025_o2_n_spl_00;
  wire n6025_o2_n_spl_1;
  wire n1003_o2_p_spl_;
  wire n1003_o2_n_spl_;
  wire g965_n_spl_;
  wire g966_p_spl_;
  wire g965_p_spl_;
  wire g966_n_spl_;
  wire g967_n_spl_;
  wire g967_p_spl_;
  wire g964_n_spl_;
  wire g969_p_spl_;
  wire g964_p_spl_;
  wire g969_n_spl_;
  wire g970_n_spl_;
  wire g970_p_spl_;
  wire g963_n_spl_;
  wire g972_p_spl_;
  wire g963_p_spl_;
  wire g972_n_spl_;
  wire g973_n_spl_;
  wire g973_p_spl_;
  wire g962_n_spl_;
  wire g975_p_spl_;
  wire g962_p_spl_;
  wire g975_n_spl_;
  wire g976_n_spl_;
  wire g976_p_spl_;
  wire g961_n_spl_;
  wire g978_p_spl_;
  wire g961_p_spl_;
  wire g978_n_spl_;
  wire g979_n_spl_;
  wire g979_p_spl_;
  wire g960_n_spl_;
  wire g981_p_spl_;
  wire g960_p_spl_;
  wire g981_n_spl_;
  wire g982_n_spl_;
  wire g982_p_spl_;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_01;
  wire G2_p_spl_1;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_000;
  wire G17_p_spl_001;
  wire G17_p_spl_01;
  wire G17_p_spl_010;
  wire G17_p_spl_011;
  wire G17_p_spl_1;
  wire G17_p_spl_10;
  wire G17_p_spl_100;
  wire G17_p_spl_101;
  wire G17_p_spl_11;
  wire G17_p_spl_110;
  wire G17_p_spl_111;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_1;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_000;
  wire G17_n_spl_001;
  wire G17_n_spl_01;
  wire G17_n_spl_010;
  wire G17_n_spl_011;
  wire G17_n_spl_1;
  wire G17_n_spl_10;
  wire G17_n_spl_100;
  wire G17_n_spl_101;
  wire G17_n_spl_11;
  wire G17_n_spl_110;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_000;
  wire G18_p_spl_001;
  wire G18_p_spl_01;
  wire G18_p_spl_010;
  wire G18_p_spl_011;
  wire G18_p_spl_1;
  wire G18_p_spl_10;
  wire G18_p_spl_100;
  wire G18_p_spl_101;
  wire G18_p_spl_11;
  wire G18_p_spl_110;
  wire G18_p_spl_111;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_000;
  wire G18_n_spl_001;
  wire G18_n_spl_01;
  wire G18_n_spl_010;
  wire G18_n_spl_011;
  wire G18_n_spl_1;
  wire G18_n_spl_10;
  wire G18_n_spl_100;
  wire G18_n_spl_101;
  wire G18_n_spl_11;
  wire G18_n_spl_110;
  wire G18_n_spl_111;
  wire g984_p_spl_;
  wire g907_p_spl_;
  wire n2758_lo_p_spl_;
  wire n2758_lo_p_spl_0;
  wire n2758_lo_p_spl_00;
  wire n2758_lo_p_spl_000;
  wire n2758_lo_p_spl_001;
  wire n2758_lo_p_spl_01;
  wire n2758_lo_p_spl_010;
  wire n2758_lo_p_spl_011;
  wire n2758_lo_p_spl_1;
  wire n2758_lo_p_spl_10;
  wire n2758_lo_p_spl_100;
  wire n2758_lo_p_spl_101;
  wire n2758_lo_p_spl_11;
  wire n2758_lo_n_spl_;
  wire n2758_lo_n_spl_0;
  wire n2758_lo_n_spl_00;
  wire n2758_lo_n_spl_000;
  wire n2758_lo_n_spl_001;
  wire n2758_lo_n_spl_01;
  wire n2758_lo_n_spl_010;
  wire n2758_lo_n_spl_011;
  wire n2758_lo_n_spl_1;
  wire n2758_lo_n_spl_10;
  wire n2758_lo_n_spl_100;
  wire n2758_lo_n_spl_101;
  wire n2758_lo_n_spl_11;
  wire g985_p_spl_;
  wire g986_p_spl_;
  wire g906_p_spl_;
  wire lo010_buf_o2_p_spl_;
  wire lo010_buf_o2_p_spl_0;
  wire lo010_buf_o2_p_spl_00;
  wire lo010_buf_o2_p_spl_1;
  wire lo010_buf_o2_n_spl_;
  wire lo010_buf_o2_n_spl_0;
  wire lo010_buf_o2_n_spl_1;
  wire n601_o2_n_spl_;
  wire n625_o2_p_spl_;
  wire n601_o2_p_spl_;
  wire n625_o2_n_spl_;
  wire g995_n_spl_;
  wire g995_p_spl_;
  wire g994_n_spl_;
  wire g997_p_spl_;
  wire g994_p_spl_;
  wire g997_n_spl_;
  wire g998_n_spl_;
  wire g998_p_spl_;
  wire g993_n_spl_;
  wire g1000_p_spl_;
  wire g993_p_spl_;
  wire g1000_n_spl_;
  wire g1001_n_spl_;
  wire g1001_p_spl_;
  wire g992_n_spl_;
  wire g1003_p_spl_;
  wire g992_p_spl_;
  wire g1003_n_spl_;
  wire g1004_n_spl_;
  wire g1004_p_spl_;
  wire g991_n_spl_;
  wire g1006_p_spl_;
  wire g991_p_spl_;
  wire g1006_n_spl_;
  wire g1007_n_spl_;
  wire g1007_p_spl_;
  wire g990_n_spl_;
  wire g1009_p_spl_;
  wire g990_p_spl_;
  wire g1009_n_spl_;
  wire g1010_n_spl_;
  wire g1010_p_spl_;
  wire g959_p_spl_;
  wire g958_n_spl_;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_000;
  wire G19_p_spl_001;
  wire G19_p_spl_01;
  wire G19_p_spl_010;
  wire G19_p_spl_011;
  wire G19_p_spl_1;
  wire G19_p_spl_10;
  wire G19_p_spl_100;
  wire G19_p_spl_101;
  wire G19_p_spl_11;
  wire G19_p_spl_110;
  wire G19_p_spl_111;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_000;
  wire G19_n_spl_001;
  wire G19_n_spl_01;
  wire G19_n_spl_010;
  wire G19_n_spl_011;
  wire G19_n_spl_1;
  wire G19_n_spl_10;
  wire G19_n_spl_100;
  wire G19_n_spl_101;
  wire G19_n_spl_11;
  wire G19_n_spl_110;
  wire G19_n_spl_111;
  wire n1811_o2_n_spl_;
  wire n1811_o2_p_spl_;
  wire n6036_o2_p_spl_;
  wire n6036_o2_p_spl_0;
  wire n6036_o2_p_spl_00;
  wire n6036_o2_p_spl_1;
  wire lo094_buf_o2_p_spl_;
  wire n6036_o2_n_spl_;
  wire n6036_o2_n_spl_0;
  wire lo094_buf_o2_n_spl_;
  wire n1889_o2_p_spl_;
  wire n1889_o2_n_spl_;
  wire g1018_n_spl_;
  wire g1019_p_spl_;
  wire g1018_p_spl_;
  wire g1019_n_spl_;
  wire g1020_n_spl_;
  wire g1020_p_spl_;
  wire g1017_n_spl_;
  wire g1022_p_spl_;
  wire g1017_p_spl_;
  wire g1022_n_spl_;
  wire n6035_o2_p_spl_;
  wire n6035_o2_p_spl_0;
  wire n6035_o2_p_spl_1;
  wire lo098_buf_o2_p_spl_;
  wire lo098_buf_o2_p_spl_0;
  wire lo098_buf_o2_p_spl_00;
  wire lo098_buf_o2_p_spl_1;
  wire n6035_o2_n_spl_;
  wire n6035_o2_n_spl_0;
  wire lo098_buf_o2_n_spl_;
  wire lo098_buf_o2_n_spl_0;
  wire lo098_buf_o2_n_spl_00;
  wire lo098_buf_o2_n_spl_1;
  wire g1023_n_spl_;
  wire g1023_p_spl_;
  wire g1024_n_spl_;
  wire g1026_p_spl_;
  wire g1024_p_spl_;
  wire g1026_n_spl_;
  wire g1027_n_spl_;
  wire g1027_p_spl_;
  wire n6037_o2_p_spl_;
  wire n6037_o2_p_spl_0;
  wire n6037_o2_p_spl_1;
  wire n6037_o2_n_spl_;
  wire n6037_o2_n_spl_0;
  wire g1030_n_spl_;
  wire g1031_n_spl_;
  wire g1030_p_spl_;
  wire g1031_p_spl_;
  wire g1032_n_spl_;
  wire g1032_p_spl_;
  wire g1029_n_spl_;
  wire g1034_p_spl_;
  wire g1029_p_spl_;
  wire g1034_n_spl_;
  wire g1035_n_spl_;
  wire g1035_p_spl_;
  wire g1028_n_spl_;
  wire g1037_p_spl_;
  wire g1028_p_spl_;
  wire g1037_n_spl_;
  wire g1038_n_spl_;
  wire g1038_p_spl_;
  wire g1039_n_spl_;
  wire g1041_p_spl_;
  wire g1039_p_spl_;
  wire g1041_n_spl_;
  wire g1042_n_spl_;
  wire g1042_p_spl_;
  wire g1045_n_spl_;
  wire g1046_n_spl_;
  wire g1045_p_spl_;
  wire g1046_p_spl_;
  wire g1047_n_spl_;
  wire g1047_p_spl_;
  wire g1044_n_spl_;
  wire g1049_p_spl_;
  wire g1044_p_spl_;
  wire g1049_n_spl_;
  wire g1050_n_spl_;
  wire g1050_p_spl_;
  wire g1043_n_spl_;
  wire g1052_p_spl_;
  wire g1043_p_spl_;
  wire g1052_n_spl_;
  wire n1631_o2_n_spl_;
  wire n1631_o2_p_spl_;
  wire n6033_o2_p_spl_;
  wire n6033_o2_p_spl_0;
  wire n6033_o2_p_spl_00;
  wire n6033_o2_p_spl_1;
  wire n6033_o2_n_spl_;
  wire n6033_o2_n_spl_0;
  wire n1725_o2_p_spl_;
  wire n1725_o2_n_spl_;
  wire g1055_n_spl_;
  wire g1056_p_spl_;
  wire g1055_p_spl_;
  wire g1056_n_spl_;
  wire g1057_n_spl_;
  wire g1057_p_spl_;
  wire g1054_n_spl_;
  wire g1059_p_spl_;
  wire g1054_p_spl_;
  wire g1059_n_spl_;
  wire n6032_o2_p_spl_;
  wire n6032_o2_p_spl_0;
  wire n6032_o2_p_spl_1;
  wire n6032_o2_n_spl_;
  wire n6032_o2_n_spl_0;
  wire g1060_n_spl_;
  wire g1060_p_spl_;
  wire g1061_n_spl_;
  wire g1063_p_spl_;
  wire g1061_p_spl_;
  wire g1063_n_spl_;
  wire g1064_n_spl_;
  wire g1064_p_spl_;
  wire n6034_o2_p_spl_;
  wire n6034_o2_p_spl_0;
  wire n6034_o2_p_spl_1;
  wire n6034_o2_n_spl_;
  wire n6034_o2_n_spl_0;
  wire g1069_n_spl_;
  wire g1070_p_spl_;
  wire g1069_p_spl_;
  wire g1070_n_spl_;
  wire g1071_n_spl_;
  wire g1071_p_spl_;
  wire g1068_n_spl_;
  wire g1073_p_spl_;
  wire g1068_p_spl_;
  wire g1073_n_spl_;
  wire g1074_n_spl_;
  wire g1074_p_spl_;
  wire g1067_n_spl_;
  wire g1076_p_spl_;
  wire g1067_p_spl_;
  wire g1076_n_spl_;
  wire g1077_n_spl_;
  wire g1077_p_spl_;
  wire g1066_n_spl_;
  wire g1079_p_spl_;
  wire g1066_p_spl_;
  wire g1079_n_spl_;
  wire g1080_n_spl_;
  wire g1080_p_spl_;
  wire g1065_n_spl_;
  wire g1082_p_spl_;
  wire g1065_p_spl_;
  wire g1082_n_spl_;
  wire g1083_n_spl_;
  wire g1083_p_spl_;
  wire g1084_n_spl_;
  wire g1086_p_spl_;
  wire g1084_p_spl_;
  wire g1086_n_spl_;
  wire g1087_n_spl_;
  wire g1087_p_spl_;
  wire g1092_n_spl_;
  wire g1094_p_spl_;
  wire g1092_p_spl_;
  wire g1094_n_spl_;
  wire g1095_n_spl_;
  wire g1095_p_spl_;
  wire g1091_n_spl_;
  wire g1097_p_spl_;
  wire g1091_p_spl_;
  wire g1097_n_spl_;
  wire g1098_n_spl_;
  wire g1098_p_spl_;
  wire g1090_n_spl_;
  wire g1100_p_spl_;
  wire g1090_p_spl_;
  wire g1100_n_spl_;
  wire g1101_n_spl_;
  wire g1101_p_spl_;
  wire g1089_n_spl_;
  wire g1103_p_spl_;
  wire g1089_p_spl_;
  wire g1103_n_spl_;
  wire g1104_n_spl_;
  wire g1104_p_spl_;
  wire g1088_n_spl_;
  wire g1106_p_spl_;
  wire g1088_p_spl_;
  wire g1106_n_spl_;
  wire n6029_o2_p_spl_;
  wire n6029_o2_p_spl_0;
  wire n6029_o2_p_spl_00;
  wire n6029_o2_p_spl_1;
  wire n6029_o2_n_spl_;
  wire n6029_o2_n_spl_0;
  wire n6029_o2_n_spl_1;
  wire n1420_o2_p_spl_;
  wire n1420_o2_n_spl_;
  wire g1108_n_spl_;
  wire g1109_p_spl_;
  wire g1108_p_spl_;
  wire g1109_n_spl_;
  wire g1110_n_spl_;
  wire g1110_p_spl_;
  wire n6030_o2_p_spl_;
  wire n6030_o2_p_spl_0;
  wire n6030_o2_p_spl_00;
  wire n6030_o2_p_spl_1;
  wire n6030_o2_n_spl_;
  wire n6030_o2_n_spl_0;
  wire n1529_o2_p_spl_;
  wire n1529_o2_n_spl_;
  wire g1112_n_spl_;
  wire g1113_p_spl_;
  wire g1112_p_spl_;
  wire g1113_n_spl_;
  wire g1114_n_spl_;
  wire g1114_p_spl_;
  wire g1111_n_spl_;
  wire g1116_p_spl_;
  wire g1111_p_spl_;
  wire g1116_n_spl_;
  wire g1117_n_spl_;
  wire g1117_p_spl_;
  wire g1118_n_spl_;
  wire g1120_p_spl_;
  wire g1118_p_spl_;
  wire g1120_n_spl_;
  wire g1121_n_spl_;
  wire g1121_p_spl_;
  wire n6031_o2_p_spl_;
  wire n6031_o2_p_spl_0;
  wire n6031_o2_p_spl_1;
  wire n6031_o2_n_spl_;
  wire n6031_o2_n_spl_0;
  wire g1126_n_spl_;
  wire g1127_p_spl_;
  wire g1126_p_spl_;
  wire g1127_n_spl_;
  wire g1128_n_spl_;
  wire g1128_p_spl_;
  wire g1125_n_spl_;
  wire g1130_p_spl_;
  wire g1125_p_spl_;
  wire g1130_n_spl_;
  wire g1131_n_spl_;
  wire g1131_p_spl_;
  wire g1124_n_spl_;
  wire g1133_p_spl_;
  wire g1124_p_spl_;
  wire g1133_n_spl_;
  wire g1134_n_spl_;
  wire g1134_p_spl_;
  wire g1123_n_spl_;
  wire g1136_p_spl_;
  wire g1123_p_spl_;
  wire g1136_n_spl_;
  wire g1137_n_spl_;
  wire g1137_p_spl_;
  wire g1122_n_spl_;
  wire g1139_p_spl_;
  wire g1122_p_spl_;
  wire g1139_n_spl_;
  wire g1140_n_spl_;
  wire g1140_p_spl_;
  wire g1141_n_spl_;
  wire g1143_p_spl_;
  wire g1141_p_spl_;
  wire g1143_n_spl_;
  wire g1144_n_spl_;
  wire g1144_p_spl_;
  wire g1149_n_spl_;
  wire g1151_p_spl_;
  wire g1149_p_spl_;
  wire g1151_n_spl_;
  wire g1152_n_spl_;
  wire g1152_p_spl_;
  wire g1148_n_spl_;
  wire g1154_p_spl_;
  wire g1148_p_spl_;
  wire g1154_n_spl_;
  wire g1155_n_spl_;
  wire g1155_p_spl_;
  wire g1147_n_spl_;
  wire g1157_p_spl_;
  wire g1147_p_spl_;
  wire g1157_n_spl_;
  wire g1158_n_spl_;
  wire g1158_p_spl_;
  wire g1146_n_spl_;
  wire g1160_p_spl_;
  wire g1146_p_spl_;
  wire g1160_n_spl_;
  wire g1161_n_spl_;
  wire g1161_p_spl_;
  wire g1145_n_spl_;
  wire g1163_p_spl_;
  wire g1145_p_spl_;
  wire g1163_n_spl_;
  wire n6026_o2_p_spl_;
  wire n6026_o2_p_spl_0;
  wire n6026_o2_p_spl_00;
  wire n6026_o2_p_spl_01;
  wire n6026_o2_p_spl_1;
  wire n6026_o2_n_spl_;
  wire n6026_o2_n_spl_0;
  wire n6026_o2_n_spl_00;
  wire n6026_o2_n_spl_1;
  wire n1097_o2_p_spl_;
  wire n1097_o2_n_spl_;
  wire g1165_n_spl_;
  wire g1166_p_spl_;
  wire g1165_p_spl_;
  wire g1166_n_spl_;
  wire g1167_n_spl_;
  wire g1167_p_spl_;
  wire n6027_o2_p_spl_;
  wire n6027_o2_p_spl_0;
  wire n6027_o2_p_spl_00;
  wire n6027_o2_p_spl_01;
  wire n6027_o2_p_spl_1;
  wire n6027_o2_n_spl_;
  wire n6027_o2_n_spl_0;
  wire n6027_o2_n_spl_1;
  wire n1199_o2_p_spl_;
  wire n1199_o2_n_spl_;
  wire g1169_n_spl_;
  wire g1170_p_spl_;
  wire g1169_p_spl_;
  wire g1170_n_spl_;
  wire g1171_n_spl_;
  wire g1171_p_spl_;
  wire g1168_n_spl_;
  wire g1173_p_spl_;
  wire g1168_p_spl_;
  wire g1173_n_spl_;
  wire g1174_n_spl_;
  wire g1174_p_spl_;
  wire g1175_n_spl_;
  wire g1177_p_spl_;
  wire g1175_p_spl_;
  wire g1177_n_spl_;
  wire g1178_n_spl_;
  wire g1178_p_spl_;
  wire n6028_o2_p_spl_;
  wire n6028_o2_p_spl_0;
  wire n6028_o2_p_spl_00;
  wire n6028_o2_p_spl_1;
  wire n6028_o2_n_spl_;
  wire n6028_o2_n_spl_0;
  wire n6028_o2_n_spl_1;
  wire n1309_o2_p_spl_;
  wire n1309_o2_n_spl_;
  wire g1182_n_spl_;
  wire g1183_p_spl_;
  wire g1182_p_spl_;
  wire g1183_n_spl_;
  wire g1184_n_spl_;
  wire g1184_p_spl_;
  wire g1181_n_spl_;
  wire g1186_p_spl_;
  wire g1181_p_spl_;
  wire g1186_n_spl_;
  wire g1187_n_spl_;
  wire g1187_p_spl_;
  wire g1180_n_spl_;
  wire g1189_p_spl_;
  wire g1180_p_spl_;
  wire g1189_n_spl_;
  wire g1190_n_spl_;
  wire g1190_p_spl_;
  wire g1179_n_spl_;
  wire g1192_p_spl_;
  wire g1179_p_spl_;
  wire g1192_n_spl_;
  wire g1193_n_spl_;
  wire g1193_p_spl_;
  wire g1194_n_spl_;
  wire g1196_p_spl_;
  wire g1194_p_spl_;
  wire g1196_n_spl_;
  wire g1197_n_spl_;
  wire g1197_p_spl_;
  wire g1202_n_spl_;
  wire g1204_p_spl_;
  wire g1202_p_spl_;
  wire g1204_n_spl_;
  wire g1205_n_spl_;
  wire g1205_p_spl_;
  wire g1201_n_spl_;
  wire g1207_p_spl_;
  wire g1201_p_spl_;
  wire g1207_n_spl_;
  wire g1208_n_spl_;
  wire g1208_p_spl_;
  wire g1200_n_spl_;
  wire g1210_p_spl_;
  wire g1200_p_spl_;
  wire g1210_n_spl_;
  wire g1211_n_spl_;
  wire g1211_p_spl_;
  wire g1199_n_spl_;
  wire g1213_p_spl_;
  wire g1199_p_spl_;
  wire g1213_n_spl_;
  wire g1214_n_spl_;
  wire g1214_p_spl_;
  wire g1198_n_spl_;
  wire g1216_p_spl_;
  wire g1198_p_spl_;
  wire g1216_n_spl_;
  wire g1217_n_spl_;
  wire g1217_p_spl_;
  wire g1218_n_spl_;
  wire g1220_p_spl_;
  wire g1218_p_spl_;
  wire g1220_n_spl_;
  wire g1221_n_spl_;
  wire g1221_p_spl_;
  wire g1226_n_spl_;
  wire g1228_p_spl_;
  wire g1226_p_spl_;
  wire g1228_n_spl_;
  wire g1229_n_spl_;
  wire g1229_p_spl_;
  wire g1225_n_spl_;
  wire g1231_p_spl_;
  wire g1225_p_spl_;
  wire g1231_n_spl_;
  wire g1232_n_spl_;
  wire g1232_p_spl_;
  wire g1224_n_spl_;
  wire g1234_p_spl_;
  wire g1224_p_spl_;
  wire g1234_n_spl_;
  wire g1235_n_spl_;
  wire g1235_p_spl_;
  wire g1223_n_spl_;
  wire g1237_p_spl_;
  wire g1223_p_spl_;
  wire g1237_n_spl_;
  wire g1238_n_spl_;
  wire g1238_p_spl_;
  wire g1222_n_spl_;
  wire g1240_p_spl_;
  wire g1222_p_spl_;
  wire g1240_n_spl_;
  wire g1012_p_spl_;
  wire g988_p_spl_;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_01;
  wire G3_p_spl_1;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_1;
  wire g1243_p_spl_;
  wire g1244_p_spl_;
  wire g1243_n_spl_;
  wire g1244_n_spl_;
  wire g1245_n_spl_;
  wire g1245_n_spl_0;
  wire g1245_p_spl_;
  wire g1245_p_spl_0;
  wire g989_n_spl_;
  wire g1247_n_spl_;
  wire g989_p_spl_;
  wire g989_p_spl_0;
  wire g1247_p_spl_;
  wire g1248_n_spl_;
  wire g1248_p_spl_;
  wire g987_p_spl_;
  wire g1257_n_spl_;
  wire g1259_p_spl_;
  wire g1257_p_spl_;
  wire g1259_n_spl_;
  wire g1260_n_spl_;
  wire g1260_p_spl_;
  wire g1256_n_spl_;
  wire g1262_p_spl_;
  wire g1256_p_spl_;
  wire g1262_n_spl_;
  wire g1263_n_spl_;
  wire g1263_p_spl_;
  wire g1255_n_spl_;
  wire g1265_p_spl_;
  wire g1255_p_spl_;
  wire g1265_n_spl_;
  wire g1266_n_spl_;
  wire g1266_p_spl_;
  wire g1254_n_spl_;
  wire g1268_p_spl_;
  wire g1254_p_spl_;
  wire g1268_n_spl_;
  wire g1269_n_spl_;
  wire g1269_p_spl_;
  wire g1253_n_spl_;
  wire g1271_p_spl_;
  wire g1253_p_spl_;
  wire g1271_n_spl_;
  wire g1272_n_spl_;
  wire g1272_p_spl_;
  wire g1252_n_spl_;
  wire g1274_p_spl_;
  wire g1252_p_spl_;
  wire g1274_n_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire n1374_o2_n_spl_;
  wire n1392_o2_p_spl_;
  wire n1374_o2_p_spl_;
  wire n1392_o2_n_spl_;
  wire g1279_n_spl_;
  wire g1279_p_spl_;
  wire n1488_o2_n_spl_;
  wire n1501_o2_p_spl_;
  wire n1488_o2_p_spl_;
  wire n1501_o2_n_spl_;
  wire g1281_n_spl_;
  wire g1281_p_spl_;
  wire g1280_n_spl_;
  wire g1283_p_spl_;
  wire g1280_p_spl_;
  wire g1283_n_spl_;
  wire lo050_buf_o2_p_spl_;
  wire lo050_buf_o2_p_spl_0;
  wire lo050_buf_o2_p_spl_1;
  wire lo050_buf_o2_n_spl_;
  wire lo050_buf_o2_n_spl_0;
  wire g1284_n_spl_;
  wire g1284_p_spl_;
  wire g1285_n_spl_;
  wire g1287_p_spl_;
  wire g1285_p_spl_;
  wire g1287_n_spl_;
  wire g1288_n_spl_;
  wire g1288_p_spl_;
  wire lo054_buf_o2_p_spl_;
  wire lo054_buf_o2_p_spl_0;
  wire lo054_buf_o2_n_spl_;
  wire lo054_buf_o2_n_spl_0;
  wire lo058_buf_o2_p_spl_;
  wire lo058_buf_o2_p_spl_0;
  wire lo058_buf_o2_p_spl_1;
  wire lo058_buf_o2_n_spl_;
  wire lo058_buf_o2_n_spl_0;
  wire n1602_o2_n_spl_;
  wire n1603_o2_n_spl_;
  wire n1602_o2_p_spl_;
  wire n1603_o2_p_spl_;
  wire g1293_n_spl_;
  wire g1293_p_spl_;
  wire g1292_n_spl_;
  wire g1295_p_spl_;
  wire g1292_p_spl_;
  wire g1295_n_spl_;
  wire g1296_n_spl_;
  wire g1296_p_spl_;
  wire g1291_n_spl_;
  wire g1298_p_spl_;
  wire g1291_p_spl_;
  wire g1298_n_spl_;
  wire g1299_n_spl_;
  wire g1299_p_spl_;
  wire g1290_n_spl_;
  wire g1301_p_spl_;
  wire g1290_p_spl_;
  wire g1301_n_spl_;
  wire g1302_n_spl_;
  wire g1302_p_spl_;
  wire g1289_n_spl_;
  wire g1304_p_spl_;
  wire g1289_p_spl_;
  wire g1304_n_spl_;
  wire g1305_n_spl_;
  wire g1305_p_spl_;
  wire g1306_n_spl_;
  wire g1308_p_spl_;
  wire g1306_p_spl_;
  wire g1308_n_spl_;
  wire g1309_n_spl_;
  wire g1309_p_spl_;
  wire lo062_buf_o2_p_spl_;
  wire lo062_buf_o2_p_spl_0;
  wire lo062_buf_o2_n_spl_;
  wire lo062_buf_o2_n_spl_0;
  wire g1314_n_spl_;
  wire g1315_n_spl_;
  wire g1314_p_spl_;
  wire g1315_p_spl_;
  wire g1316_n_spl_;
  wire g1316_p_spl_;
  wire g1313_n_spl_;
  wire g1318_p_spl_;
  wire g1313_p_spl_;
  wire g1318_n_spl_;
  wire g1319_n_spl_;
  wire g1319_p_spl_;
  wire g1312_n_spl_;
  wire g1321_p_spl_;
  wire g1312_p_spl_;
  wire g1321_n_spl_;
  wire g1322_n_spl_;
  wire g1322_p_spl_;
  wire g1311_n_spl_;
  wire g1324_p_spl_;
  wire g1311_p_spl_;
  wire g1324_n_spl_;
  wire g1325_n_spl_;
  wire g1325_p_spl_;
  wire g1310_n_spl_;
  wire g1327_p_spl_;
  wire g1310_p_spl_;
  wire g1327_n_spl_;
  wire n1045_o2_n_spl_;
  wire n1069_o2_p_spl_;
  wire n1045_o2_p_spl_;
  wire n1069_o2_n_spl_;
  wire g1329_n_spl_;
  wire g1329_p_spl_;
  wire n1147_o2_n_spl_;
  wire n1171_o2_p_spl_;
  wire n1147_o2_p_spl_;
  wire n1171_o2_n_spl_;
  wire g1331_n_spl_;
  wire g1331_p_spl_;
  wire g1330_n_spl_;
  wire g1333_p_spl_;
  wire g1330_p_spl_;
  wire g1333_n_spl_;
  wire lo038_buf_o2_p_spl_;
  wire lo038_buf_o2_p_spl_0;
  wire lo038_buf_o2_p_spl_00;
  wire lo038_buf_o2_p_spl_1;
  wire lo038_buf_o2_n_spl_;
  wire lo038_buf_o2_n_spl_0;
  wire lo038_buf_o2_n_spl_1;
  wire g1334_n_spl_;
  wire g1334_p_spl_;
  wire g1335_n_spl_;
  wire g1337_p_spl_;
  wire g1335_p_spl_;
  wire g1337_n_spl_;
  wire g1338_n_spl_;
  wire g1338_p_spl_;
  wire lo042_buf_o2_p_spl_;
  wire lo042_buf_o2_p_spl_0;
  wire lo042_buf_o2_p_spl_1;
  wire lo042_buf_o2_n_spl_;
  wire lo042_buf_o2_n_spl_0;
  wire lo042_buf_o2_n_spl_1;
  wire n1257_o2_n_spl_;
  wire n1281_o2_p_spl_;
  wire n1257_o2_p_spl_;
  wire n1281_o2_n_spl_;
  wire g1342_n_spl_;
  wire g1342_p_spl_;
  wire g1341_n_spl_;
  wire g1344_p_spl_;
  wire g1341_p_spl_;
  wire g1344_n_spl_;
  wire g1345_n_spl_;
  wire g1345_p_spl_;
  wire g1340_n_spl_;
  wire g1347_p_spl_;
  wire g1340_p_spl_;
  wire g1347_n_spl_;
  wire g1348_n_spl_;
  wire g1348_p_spl_;
  wire g1339_n_spl_;
  wire g1350_p_spl_;
  wire g1339_p_spl_;
  wire g1350_n_spl_;
  wire g1351_n_spl_;
  wire g1351_p_spl_;
  wire g1352_n_spl_;
  wire g1354_p_spl_;
  wire g1352_p_spl_;
  wire g1354_n_spl_;
  wire g1355_n_spl_;
  wire g1355_p_spl_;
  wire lo046_buf_o2_p_spl_;
  wire lo046_buf_o2_p_spl_0;
  wire lo046_buf_o2_p_spl_1;
  wire lo046_buf_o2_n_spl_;
  wire lo046_buf_o2_n_spl_0;
  wire g1360_n_spl_;
  wire g1362_p_spl_;
  wire g1360_p_spl_;
  wire g1362_n_spl_;
  wire g1363_n_spl_;
  wire g1363_p_spl_;
  wire g1359_n_spl_;
  wire g1365_p_spl_;
  wire g1359_p_spl_;
  wire g1365_n_spl_;
  wire g1366_n_spl_;
  wire g1366_p_spl_;
  wire g1358_n_spl_;
  wire g1368_p_spl_;
  wire g1358_p_spl_;
  wire g1368_n_spl_;
  wire g1369_n_spl_;
  wire g1369_p_spl_;
  wire g1357_n_spl_;
  wire g1371_p_spl_;
  wire g1357_p_spl_;
  wire g1371_n_spl_;
  wire g1372_n_spl_;
  wire g1372_p_spl_;
  wire g1356_n_spl_;
  wire g1374_p_spl_;
  wire g1356_p_spl_;
  wire g1374_n_spl_;
  wire g1375_n_spl_;
  wire g1375_p_spl_;
  wire g1376_n_spl_;
  wire g1378_p_spl_;
  wire g1376_p_spl_;
  wire g1378_n_spl_;
  wire g1379_n_spl_;
  wire g1379_p_spl_;
  wire g1384_n_spl_;
  wire g1386_p_spl_;
  wire g1384_p_spl_;
  wire g1386_n_spl_;
  wire g1387_n_spl_;
  wire g1387_p_spl_;
  wire g1383_n_spl_;
  wire g1389_p_spl_;
  wire g1383_p_spl_;
  wire g1389_n_spl_;
  wire g1390_n_spl_;
  wire g1390_p_spl_;
  wire g1382_n_spl_;
  wire g1392_p_spl_;
  wire g1382_p_spl_;
  wire g1392_n_spl_;
  wire g1393_n_spl_;
  wire g1393_p_spl_;
  wire g1381_n_spl_;
  wire g1395_p_spl_;
  wire g1381_p_spl_;
  wire g1395_n_spl_;
  wire g1396_n_spl_;
  wire g1396_p_spl_;
  wire g1380_n_spl_;
  wire g1398_p_spl_;
  wire g1380_p_spl_;
  wire g1398_n_spl_;
  wire g1250_p_spl_;
  wire g1016_p_spl_;
  wire n2833_lo_n_spl_;
  wire n2833_lo_n_spl_0;
  wire n2833_lo_n_spl_00;
  wire n2833_lo_n_spl_1;
  wire n2770_lo_n_spl_;
  wire n2770_lo_n_spl_0;
  wire n2770_lo_n_spl_00;
  wire n2770_lo_n_spl_000;
  wire n2770_lo_n_spl_001;
  wire n2770_lo_n_spl_01;
  wire n2770_lo_n_spl_010;
  wire n2770_lo_n_spl_1;
  wire n2770_lo_n_spl_10;
  wire n2770_lo_n_spl_11;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_000;
  wire G20_n_spl_001;
  wire G20_n_spl_01;
  wire G20_n_spl_010;
  wire G20_n_spl_011;
  wire G20_n_spl_1;
  wire G20_n_spl_10;
  wire G20_n_spl_100;
  wire G20_n_spl_101;
  wire G20_n_spl_11;
  wire G20_n_spl_110;
  wire g946_n_spl_;
  wire g1404_n_spl_;
  wire g1406_p_spl_;
  wire g934_n_spl_;
  wire g1409_n_spl_;
  wire g1411_p_spl_;
  wire g922_n_spl_;
  wire g1414_n_spl_;
  wire g1416_p_spl_;
  wire g919_n_spl_;
  wire g1419_n_spl_;
  wire g1421_p_spl_;
  wire g915_n_spl_;
  wire g1424_n_spl_;
  wire g1426_p_spl_;
  wire g911_n_spl_;
  wire g1429_n_spl_;
  wire g1431_p_spl_;
  wire g1013_n_spl_;
  wire g1015_p_spl_;
  wire n2833_lo_p_spl_;
  wire n2833_lo_p_spl_0;
  wire n2833_lo_p_spl_00;
  wire n2833_lo_p_spl_1;
  wire g1241_n_spl_;
  wire g1164_n_spl_;
  wire g1107_n_spl_;
  wire g1053_n_spl_;
  wire g1459_n_spl_;
  wire g1461_p_spl_;
  wire g1459_p_spl_;
  wire g1461_n_spl_;
  wire g1462_n_spl_;
  wire g1462_p_spl_;
  wire g1458_n_spl_;
  wire g1464_p_spl_;
  wire g1458_p_spl_;
  wire g1464_n_spl_;
  wire g1465_n_spl_;
  wire g1465_p_spl_;
  wire g1457_n_spl_;
  wire g1467_p_spl_;
  wire g1457_p_spl_;
  wire g1467_n_spl_;
  wire g1468_n_spl_;
  wire g1468_p_spl_;
  wire g1456_n_spl_;
  wire g1470_p_spl_;
  wire g1456_p_spl_;
  wire g1470_n_spl_;
  wire g1471_n_spl_;
  wire g1471_p_spl_;
  wire g1455_n_spl_;
  wire g1473_p_spl_;
  wire g1454_n_spl_;
  wire g1476_p_spl_;
  wire g1480_n_spl_;
  wire g1482_p_spl_;
  wire g1480_p_spl_;
  wire g1482_n_spl_;
  wire g1483_n_spl_;
  wire g1479_n_spl_;
  wire g1485_p_spl_;
  wire g1479_p_spl_;
  wire g1485_n_spl_;
  wire g1486_n_spl_;
  wire g1492_n_spl_;
  wire g1494_p_spl_;
  wire g1492_p_spl_;
  wire g1494_n_spl_;
  wire g1495_n_spl_;
  wire g1491_n_spl_;
  wire g1497_p_spl_;
  wire g1491_p_spl_;
  wire g1497_n_spl_;
  wire g1498_n_spl_;
  wire g1504_n_spl_;
  wire g1506_p_spl_;
  wire g1504_p_spl_;
  wire g1506_n_spl_;
  wire g1507_n_spl_;
  wire g1503_n_spl_;
  wire g1509_p_spl_;
  wire g1503_p_spl_;
  wire g1509_n_spl_;
  wire g1510_n_spl_;
  wire g1278_n_spl_;
  wire n2770_lo_p_spl_;
  wire n2770_lo_p_spl_0;
  wire n2770_lo_p_spl_00;
  wire n2770_lo_p_spl_000;
  wire n2770_lo_p_spl_001;
  wire n2770_lo_p_spl_01;
  wire n2770_lo_p_spl_1;
  wire n2770_lo_p_spl_10;
  wire n2770_lo_p_spl_11;
  wire g1399_n_spl_;
  wire g1328_n_spl_;
  wire g1526_n_spl_;
  wire g1527_n_spl_;
  wire g1526_p_spl_;
  wire g1527_p_spl_;
  wire g1528_p_spl_;
  wire g1525_n_spl_;
  wire g1530_p_spl_;
  wire g1525_p_spl_;
  wire g1530_n_spl_;
  wire g1531_p_spl_;
  wire g1537_n_spl_;
  wire g1539_p_spl_;
  wire g1537_p_spl_;
  wire g1539_n_spl_;
  wire g1540_p_spl_;
  wire g1536_n_spl_;
  wire g1542_p_spl_;
  wire g1536_p_spl_;
  wire g1542_n_spl_;
  wire g1543_p_spl_;
  wire g1242_p_spl_;
  wire lo014_buf_o2_p_spl_;
  wire lo014_buf_o2_p_spl_0;
  wire lo014_buf_o2_p_spl_00;
  wire lo014_buf_o2_p_spl_1;
  wire lo014_buf_o2_n_spl_;
  wire lo014_buf_o2_n_spl_0;
  wire lo014_buf_o2_n_spl_1;
  wire n655_o2_n_spl_;
  wire n679_o2_p_spl_;
  wire n655_o2_p_spl_;
  wire n679_o2_n_spl_;
  wire g1554_n_spl_;
  wire g1554_p_spl_;
  wire g1553_n_spl_;
  wire g1556_p_spl_;
  wire g1553_p_spl_;
  wire g1556_n_spl_;
  wire g1557_n_spl_;
  wire g1557_p_spl_;
  wire g1552_n_spl_;
  wire g1559_p_spl_;
  wire g1552_p_spl_;
  wire g1559_n_spl_;
  wire g1560_n_spl_;
  wire g1560_p_spl_;
  wire g1551_n_spl_;
  wire g1562_p_spl_;
  wire g1551_p_spl_;
  wire g1562_n_spl_;
  wire g1563_n_spl_;
  wire g1563_p_spl_;
  wire g1550_n_spl_;
  wire g1565_p_spl_;
  wire g1550_p_spl_;
  wire g1565_n_spl_;
  wire g1566_n_spl_;
  wire g1566_p_spl_;
  wire g1549_n_spl_;
  wire g1568_p_spl_;
  wire g1549_p_spl_;
  wire g1568_n_spl_;
  wire g1569_n_spl_;
  wire g1569_p_spl_;
  wire g1548_n_spl_;
  wire g1571_p_spl_;
  wire g1548_p_spl_;
  wire g1571_n_spl_;
  wire g1572_n_spl_;
  wire g1572_p_spl_;
  wire g1547_n_spl_;
  wire g1574_p_spl_;
  wire g1400_p_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_1;
  wire g1580_p_spl_;
  wire g1581_p_spl_;
  wire g1580_n_spl_;
  wire g1581_n_spl_;
  wire g1582_n_spl_;
  wire g1582_n_spl_0;
  wire g1582_p_spl_;
  wire g1582_p_spl_0;
  wire g1584_n_spl_;
  wire g1584_p_spl_;
  wire g1585_n_spl_;
  wire g1585_p_spl_;
  wire g1579_n_spl_;
  wire g1587_p_spl_;
  wire g1579_p_spl_;
  wire g1587_n_spl_;
  wire g1588_n_spl_;
  wire g1588_p_spl_;
  wire g1578_n_spl_;
  wire g1590_p_spl_;
  wire g1603_n_spl_;
  wire g1605_p_spl_;
  wire g1603_p_spl_;
  wire g1605_n_spl_;
  wire g1606_n_spl_;
  wire g1606_p_spl_;
  wire g1602_n_spl_;
  wire g1608_p_spl_;
  wire g1602_p_spl_;
  wire g1608_n_spl_;
  wire g1609_n_spl_;
  wire g1609_p_spl_;
  wire g1601_n_spl_;
  wire g1611_p_spl_;
  wire g1601_p_spl_;
  wire g1611_n_spl_;
  wire g1612_n_spl_;
  wire g1616_n_spl_;
  wire g1618_n_spl_;
  wire g1620_p_spl_;
  wire g1618_p_spl_;
  wire g1620_n_spl_;
  wire g1621_n_spl_;
  wire g1625_n_spl_;
  wire g1477_p_spl_;
  wire g1401_n_spl_;
  wire g1515_p_spl_;
  wire g1402_n_spl_;
  wire g1577_p_spl_;
  wire g1403_n_spl_;
  wire g1593_p_spl_;
  wire g1438_n_spl_;
  wire g1442_n_spl_;
  wire g1446_n_spl_;
  wire g1450_n_spl_;
  wire g1453_n_spl_;
  wire g1489_n_spl_;
  wire g1501_n_spl_;
  wire g1513_n_spl_;
  wire g1630_p_spl_;
  wire lo018_buf_o2_p_spl_;
  wire lo018_buf_o2_p_spl_0;
  wire lo018_buf_o2_p_spl_00;
  wire lo018_buf_o2_p_spl_1;
  wire lo018_buf_o2_n_spl_;
  wire lo018_buf_o2_n_spl_0;
  wire lo018_buf_o2_n_spl_1;
  wire n717_o2_n_spl_;
  wire n741_o2_p_spl_;
  wire n717_o2_p_spl_;
  wire n741_o2_n_spl_;
  wire g1661_n_spl_;
  wire g1661_p_spl_;
  wire g1660_n_spl_;
  wire g1663_p_spl_;
  wire g1660_p_spl_;
  wire g1663_n_spl_;
  wire g1664_n_spl_;
  wire g1664_p_spl_;
  wire g1659_n_spl_;
  wire g1666_p_spl_;
  wire g1659_p_spl_;
  wire g1666_n_spl_;
  wire g1667_n_spl_;
  wire g1667_p_spl_;
  wire g1658_n_spl_;
  wire g1669_p_spl_;
  wire g1658_p_spl_;
  wire g1669_n_spl_;
  wire g1670_n_spl_;
  wire g1670_p_spl_;
  wire g1657_n_spl_;
  wire g1672_p_spl_;
  wire g1657_p_spl_;
  wire g1672_n_spl_;
  wire g1673_n_spl_;
  wire g1673_p_spl_;
  wire g1656_n_spl_;
  wire g1675_p_spl_;
  wire g1656_p_spl_;
  wire g1675_n_spl_;
  wire g1676_n_spl_;
  wire g1676_p_spl_;
  wire g1655_n_spl_;
  wire g1678_p_spl_;
  wire g1655_p_spl_;
  wire g1678_n_spl_;
  wire g1679_n_spl_;
  wire g1679_p_spl_;
  wire g1654_n_spl_;
  wire g1681_p_spl_;
  wire g1654_p_spl_;
  wire g1681_n_spl_;
  wire g1682_n_spl_;
  wire g1685_n_spl_;
  wire g1546_n_spl_;
  wire g1688_n_spl_;
  wire g1690_p_spl_;
  wire g1534_n_spl_;
  wire g1693_n_spl_;
  wire g1695_p_spl_;
  wire g1698_n_spl_;
  wire g1699_n_spl_;
  wire g1523_n_spl_;
  wire g1702_n_spl_;
  wire g1704_p_spl_;
  wire lo022_buf_o2_p_spl_;
  wire lo022_buf_o2_p_spl_0;
  wire lo022_buf_o2_p_spl_00;
  wire lo022_buf_o2_p_spl_1;
  wire lo022_buf_o2_n_spl_;
  wire lo022_buf_o2_n_spl_0;
  wire lo022_buf_o2_n_spl_1;
  wire n787_o2_n_spl_;
  wire n811_o2_p_spl_;
  wire n787_o2_p_spl_;
  wire n811_o2_n_spl_;
  wire g1714_n_spl_;
  wire g1714_p_spl_;
  wire g1713_n_spl_;
  wire g1716_p_spl_;
  wire g1713_p_spl_;
  wire g1716_n_spl_;
  wire g1717_n_spl_;
  wire g1717_p_spl_;
  wire g1712_n_spl_;
  wire g1719_p_spl_;
  wire g1712_p_spl_;
  wire g1719_n_spl_;
  wire g1720_n_spl_;
  wire g1720_p_spl_;
  wire g1711_n_spl_;
  wire g1722_p_spl_;
  wire g1711_p_spl_;
  wire g1722_n_spl_;
  wire g1723_n_spl_;
  wire g1723_p_spl_;
  wire g1710_n_spl_;
  wire g1725_p_spl_;
  wire g1710_p_spl_;
  wire g1725_n_spl_;
  wire g1726_n_spl_;
  wire g1726_p_spl_;
  wire g1709_n_spl_;
  wire g1728_p_spl_;
  wire g1709_p_spl_;
  wire g1728_n_spl_;
  wire g1729_n_spl_;
  wire g1729_p_spl_;
  wire g1708_n_spl_;
  wire g1731_p_spl_;
  wire g1708_p_spl_;
  wire g1731_n_spl_;
  wire g1732_n_spl_;
  wire g1732_p_spl_;
  wire g1707_n_spl_;
  wire g1734_p_spl_;
  wire g1707_p_spl_;
  wire g1734_n_spl_;
  wire g1735_p_spl_;
  wire g1739_p_spl_;
  wire lo026_buf_o2_p_spl_;
  wire lo026_buf_o2_p_spl_0;
  wire lo026_buf_o2_p_spl_00;
  wire lo026_buf_o2_p_spl_1;
  wire lo026_buf_o2_n_spl_;
  wire lo026_buf_o2_n_spl_0;
  wire lo026_buf_o2_n_spl_1;
  wire n865_o2_n_spl_;
  wire n889_o2_p_spl_;
  wire n865_o2_p_spl_;
  wire n889_o2_n_spl_;
  wire g1749_n_spl_;
  wire g1749_p_spl_;
  wire g1748_n_spl_;
  wire g1751_p_spl_;
  wire g1748_p_spl_;
  wire g1751_n_spl_;
  wire g1752_n_spl_;
  wire g1752_p_spl_;
  wire g1747_n_spl_;
  wire g1754_p_spl_;
  wire g1747_p_spl_;
  wire g1754_n_spl_;
  wire g1755_n_spl_;
  wire g1755_p_spl_;
  wire g1746_n_spl_;
  wire g1757_p_spl_;
  wire g1746_p_spl_;
  wire g1757_n_spl_;
  wire g1758_n_spl_;
  wire g1758_p_spl_;
  wire g1745_n_spl_;
  wire g1760_p_spl_;
  wire g1745_p_spl_;
  wire g1760_n_spl_;
  wire g1761_n_spl_;
  wire g1761_p_spl_;
  wire g1744_n_spl_;
  wire g1763_p_spl_;
  wire g1744_p_spl_;
  wire g1763_n_spl_;
  wire g1764_n_spl_;
  wire g1764_p_spl_;
  wire g1743_n_spl_;
  wire g1766_p_spl_;
  wire g1743_p_spl_;
  wire g1766_n_spl_;
  wire g1767_n_spl_;
  wire g1767_p_spl_;
  wire g1742_n_spl_;
  wire g1769_p_spl_;
  wire g1742_p_spl_;
  wire g1769_n_spl_;
  wire g1770_p_spl_;
  wire g1741_n_spl_;
  wire g1772_p_spl_;
  wire g1740_n_spl_;
  wire g1775_p_spl_;
  wire lo030_buf_o2_p_spl_;
  wire lo030_buf_o2_p_spl_0;
  wire lo030_buf_o2_p_spl_00;
  wire lo030_buf_o2_p_spl_1;
  wire lo030_buf_o2_n_spl_;
  wire lo030_buf_o2_n_spl_0;
  wire lo030_buf_o2_n_spl_1;
  wire n951_o2_n_spl_;
  wire n975_o2_p_spl_;
  wire n951_o2_p_spl_;
  wire n975_o2_n_spl_;
  wire g1787_n_spl_;
  wire g1787_p_spl_;
  wire g1786_n_spl_;
  wire g1789_p_spl_;
  wire g1786_p_spl_;
  wire g1789_n_spl_;
  wire g1790_n_spl_;
  wire g1790_p_spl_;
  wire g1785_n_spl_;
  wire g1792_p_spl_;
  wire g1785_p_spl_;
  wire g1792_n_spl_;
  wire g1793_n_spl_;
  wire g1793_p_spl_;
  wire g1784_n_spl_;
  wire g1795_p_spl_;
  wire g1784_p_spl_;
  wire g1795_n_spl_;
  wire g1796_n_spl_;
  wire g1796_p_spl_;
  wire g1783_n_spl_;
  wire g1798_p_spl_;
  wire g1783_p_spl_;
  wire g1798_n_spl_;
  wire g1799_n_spl_;
  wire g1799_p_spl_;
  wire g1782_n_spl_;
  wire g1801_p_spl_;
  wire g1782_p_spl_;
  wire g1801_n_spl_;
  wire g1802_n_spl_;
  wire g1802_p_spl_;
  wire g1781_n_spl_;
  wire g1804_p_spl_;
  wire g1781_p_spl_;
  wire g1804_n_spl_;
  wire g1805_n_spl_;
  wire g1805_p_spl_;
  wire g1780_n_spl_;
  wire g1807_p_spl_;
  wire g1780_p_spl_;
  wire g1807_n_spl_;
  wire g1808_p_spl_;
  wire g1779_n_spl_;
  wire g1810_p_spl_;
  wire g1778_n_spl_;
  wire g1813_p_spl_;
  wire lo034_buf_o2_p_spl_;
  wire lo034_buf_o2_p_spl_0;
  wire lo034_buf_o2_p_spl_00;
  wire lo034_buf_o2_p_spl_1;
  wire lo034_buf_o2_n_spl_;
  wire lo034_buf_o2_n_spl_0;
  wire lo034_buf_o2_n_spl_1;
  wire g1824_n_spl_;
  wire g1826_p_spl_;
  wire g1824_p_spl_;
  wire g1826_n_spl_;
  wire g1827_n_spl_;
  wire g1827_p_spl_;
  wire g1823_n_spl_;
  wire g1829_p_spl_;
  wire g1823_p_spl_;
  wire g1829_n_spl_;
  wire g1830_n_spl_;
  wire g1830_p_spl_;
  wire g1822_n_spl_;
  wire g1832_p_spl_;
  wire g1822_p_spl_;
  wire g1832_n_spl_;
  wire g1833_n_spl_;
  wire g1833_p_spl_;
  wire g1821_n_spl_;
  wire g1835_p_spl_;
  wire g1821_p_spl_;
  wire g1835_n_spl_;
  wire g1836_n_spl_;
  wire g1836_p_spl_;
  wire g1820_n_spl_;
  wire g1838_p_spl_;
  wire g1820_p_spl_;
  wire g1838_n_spl_;
  wire g1839_n_spl_;
  wire g1839_p_spl_;
  wire g1819_n_spl_;
  wire g1841_p_spl_;
  wire g1819_p_spl_;
  wire g1841_n_spl_;
  wire g1842_n_spl_;
  wire g1842_p_spl_;
  wire g1818_n_spl_;
  wire g1844_p_spl_;
  wire g1818_p_spl_;
  wire g1844_n_spl_;
  wire g1845_p_spl_;
  wire g1817_n_spl_;
  wire g1847_p_spl_;
  wire g1816_n_spl_;
  wire g1850_p_spl_;
  wire g1859_n_spl_;
  wire g1861_p_spl_;
  wire g1859_p_spl_;
  wire g1861_n_spl_;
  wire g1862_n_spl_;
  wire g1862_p_spl_;
  wire g1858_n_spl_;
  wire g1864_p_spl_;
  wire g1858_p_spl_;
  wire g1864_n_spl_;
  wire g1865_n_spl_;
  wire g1865_p_spl_;
  wire g1857_n_spl_;
  wire g1867_p_spl_;
  wire g1857_p_spl_;
  wire g1867_n_spl_;
  wire g1868_n_spl_;
  wire g1868_p_spl_;
  wire g1856_n_spl_;
  wire g1870_p_spl_;
  wire g1856_p_spl_;
  wire g1870_n_spl_;
  wire g1871_n_spl_;
  wire g1871_p_spl_;
  wire g1855_n_spl_;
  wire g1873_p_spl_;
  wire g1855_p_spl_;
  wire g1873_n_spl_;
  wire g1874_p_spl_;
  wire g1854_n_spl_;
  wire g1876_p_spl_;
  wire g1853_n_spl_;
  wire g1879_p_spl_;
  wire g1886_n_spl_;
  wire g1888_p_spl_;
  wire g1886_p_spl_;
  wire g1888_n_spl_;
  wire g1889_n_spl_;
  wire g1889_p_spl_;
  wire g1885_n_spl_;
  wire g1891_p_spl_;
  wire g1885_p_spl_;
  wire g1891_n_spl_;
  wire g1892_n_spl_;
  wire g1892_p_spl_;
  wire g1884_n_spl_;
  wire g1894_p_spl_;
  wire g1884_p_spl_;
  wire g1894_n_spl_;
  wire g1895_p_spl_;
  wire g1883_n_spl_;
  wire g1897_p_spl_;
  wire g1882_n_spl_;
  wire g1900_p_spl_;
  wire g1905_n_spl_;
  wire g1907_p_spl_;
  wire g1905_p_spl_;
  wire g1907_n_spl_;
  wire g1908_p_spl_;
  wire g1904_n_spl_;
  wire g1910_p_spl_;
  wire g1903_n_spl_;
  wire g1913_p_spl_;
  wire g1519_n_spl_;
  wire g1916_n_spl_;
  wire g1918_p_spl_;
  wire g1921_p_spl_;
  wire g1923_n_spl_;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_01;
  wire G5_p_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_1;
  wire g1926_p_spl_;
  wire g1927_p_spl_;
  wire g1926_n_spl_;
  wire g1927_n_spl_;
  wire g1928_n_spl_;
  wire g1928_n_spl_0;
  wire g1928_p_spl_;
  wire g1928_p_spl_0;
  wire g1930_n_spl_;
  wire g1930_p_spl_;
  wire g1931_n_spl_;
  wire g1931_p_spl_;
  wire g1932_n_spl_;
  wire g1934_p_spl_;
  wire g1932_p_spl_;
  wire g1934_n_spl_;
  wire g1935_n_spl_;
  wire g1935_p_spl_;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_01;
  wire G6_p_spl_1;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_1;
  wire g1938_p_spl_;
  wire g1939_p_spl_;
  wire g1938_n_spl_;
  wire g1939_n_spl_;
  wire g1940_n_spl_;
  wire g1940_n_spl_0;
  wire g1940_p_spl_;
  wire g1940_p_spl_0;
  wire g1942_n_spl_;
  wire g1942_p_spl_;
  wire g1943_n_spl_;
  wire g1943_p_spl_;
  wire g1937_n_spl_;
  wire g1945_p_spl_;
  wire g1937_p_spl_;
  wire g1945_n_spl_;
  wire g1946_n_spl_;
  wire g1946_p_spl_;
  wire g1936_n_spl_;
  wire g1948_p_spl_;
  wire g1936_p_spl_;
  wire g1948_n_spl_;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_000;
  wire G20_p_spl_001;
  wire G20_p_spl_01;
  wire G20_p_spl_010;
  wire G20_p_spl_011;
  wire G20_p_spl_1;
  wire G20_p_spl_10;
  wire G20_p_spl_100;
  wire G20_p_spl_101;
  wire G20_p_spl_11;
  wire G20_p_spl_110;
  wire g1949_n_spl_;
  wire g1949_p_spl_;
  wire g1950_n_spl_;
  wire g1952_p_spl_;
  wire g1950_p_spl_;
  wire g1952_n_spl_;
  wire g1953_n_spl_;
  wire g1953_p_spl_;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_01;
  wire G7_p_spl_1;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_1;
  wire g1958_p_spl_;
  wire g1959_p_spl_;
  wire g1958_n_spl_;
  wire g1959_n_spl_;
  wire g1960_n_spl_;
  wire g1960_n_spl_0;
  wire g1960_p_spl_;
  wire g1960_p_spl_0;
  wire g1962_n_spl_;
  wire g1962_p_spl_;
  wire g1963_n_spl_;
  wire g1963_p_spl_;
  wire g1957_n_spl_;
  wire g1965_p_spl_;
  wire g1957_p_spl_;
  wire g1965_n_spl_;
  wire g1966_n_spl_;
  wire g1966_p_spl_;
  wire g1956_n_spl_;
  wire g1968_p_spl_;
  wire g1956_p_spl_;
  wire g1968_n_spl_;
  wire g1969_n_spl_;
  wire g1969_p_spl_;
  wire g1955_n_spl_;
  wire g1971_p_spl_;
  wire g1955_p_spl_;
  wire g1971_n_spl_;
  wire g1972_n_spl_;
  wire g1972_p_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_01;
  wire G8_p_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_1;
  wire g1980_p_spl_;
  wire g1981_p_spl_;
  wire g1980_n_spl_;
  wire g1981_n_spl_;
  wire g1982_n_spl_;
  wire g1982_n_spl_0;
  wire g1982_p_spl_;
  wire g1982_p_spl_0;
  wire g1984_n_spl_;
  wire g1984_p_spl_;
  wire g1985_n_spl_;
  wire g1985_p_spl_;
  wire g1979_n_spl_;
  wire g1987_p_spl_;
  wire g1979_p_spl_;
  wire g1987_n_spl_;
  wire g1988_n_spl_;
  wire g1988_p_spl_;
  wire g1978_n_spl_;
  wire g1990_p_spl_;
  wire g1978_p_spl_;
  wire g1990_n_spl_;
  wire g1991_n_spl_;
  wire g1991_p_spl_;
  wire g1977_n_spl_;
  wire g1993_p_spl_;
  wire g1977_p_spl_;
  wire g1993_n_spl_;
  wire g1994_n_spl_;
  wire g1994_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_01;
  wire G9_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_1;
  wire g2002_p_spl_;
  wire g2003_p_spl_;
  wire g2002_n_spl_;
  wire g2003_n_spl_;
  wire g2004_n_spl_;
  wire g2004_n_spl_0;
  wire g2004_p_spl_;
  wire g2004_p_spl_0;
  wire g2006_n_spl_;
  wire g2006_p_spl_;
  wire g2007_n_spl_;
  wire g2007_p_spl_;
  wire g2001_n_spl_;
  wire g2009_p_spl_;
  wire g2001_p_spl_;
  wire g2009_n_spl_;
  wire g2010_n_spl_;
  wire g2010_p_spl_;
  wire g2000_n_spl_;
  wire g2012_p_spl_;
  wire g2000_p_spl_;
  wire g2012_n_spl_;
  wire g2013_n_spl_;
  wire g2013_p_spl_;
  wire g1999_n_spl_;
  wire g2015_p_spl_;
  wire g1999_p_spl_;
  wire g2015_n_spl_;
  wire g2016_n_spl_;
  wire g2016_p_spl_;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_01;
  wire G10_p_spl_1;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_1;
  wire g2024_p_spl_;
  wire g2025_p_spl_;
  wire g2024_n_spl_;
  wire g2025_n_spl_;
  wire g2026_n_spl_;
  wire g2026_n_spl_0;
  wire g2026_p_spl_;
  wire g2026_p_spl_0;
  wire g2028_n_spl_;
  wire g2028_p_spl_;
  wire g2029_n_spl_;
  wire g2029_p_spl_;
  wire g2023_n_spl_;
  wire g2031_p_spl_;
  wire g2023_p_spl_;
  wire g2031_n_spl_;
  wire g2032_n_spl_;
  wire g2032_p_spl_;
  wire g2022_n_spl_;
  wire g2034_p_spl_;
  wire g2022_p_spl_;
  wire g2034_n_spl_;
  wire g2035_n_spl_;
  wire g2035_p_spl_;
  wire g2021_n_spl_;
  wire g2037_p_spl_;
  wire g2021_p_spl_;
  wire g2037_n_spl_;
  wire g2038_n_spl_;
  wire g2038_p_spl_;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_01;
  wire G11_p_spl_1;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_1;
  wire g2046_p_spl_;
  wire g2047_p_spl_;
  wire g2046_n_spl_;
  wire g2047_n_spl_;
  wire g2048_n_spl_;
  wire g2048_n_spl_0;
  wire g2048_p_spl_;
  wire g2048_p_spl_0;
  wire g2050_n_spl_;
  wire g2050_p_spl_;
  wire g2051_n_spl_;
  wire g2051_p_spl_;
  wire g2045_n_spl_;
  wire g2053_p_spl_;
  wire g2045_p_spl_;
  wire g2053_n_spl_;
  wire g2054_n_spl_;
  wire g2054_p_spl_;
  wire g2044_n_spl_;
  wire g2056_p_spl_;
  wire g2044_p_spl_;
  wire g2056_n_spl_;
  wire g2057_n_spl_;
  wire g2057_p_spl_;
  wire g2043_n_spl_;
  wire g2059_p_spl_;
  wire g2043_p_spl_;
  wire g2059_n_spl_;
  wire g2060_n_spl_;
  wire g2060_p_spl_;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_01;
  wire G12_p_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_1;
  wire g2068_p_spl_;
  wire g2069_p_spl_;
  wire g2068_n_spl_;
  wire g2069_n_spl_;
  wire g2070_n_spl_;
  wire g2070_n_spl_0;
  wire g2070_p_spl_;
  wire g2070_p_spl_0;
  wire g2072_n_spl_;
  wire g2072_p_spl_;
  wire g2073_n_spl_;
  wire g2073_p_spl_;
  wire g2067_n_spl_;
  wire g2075_p_spl_;
  wire g2067_p_spl_;
  wire g2075_n_spl_;
  wire g2076_n_spl_;
  wire g2076_p_spl_;
  wire g2066_n_spl_;
  wire g2078_p_spl_;
  wire g2066_p_spl_;
  wire g2078_n_spl_;
  wire g2079_n_spl_;
  wire g2079_p_spl_;
  wire g2065_n_spl_;
  wire g2081_p_spl_;
  wire g2065_p_spl_;
  wire g2081_n_spl_;
  wire g2082_n_spl_;
  wire g2082_p_spl_;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_01;
  wire G13_p_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_1;
  wire g2090_p_spl_;
  wire g2091_p_spl_;
  wire g2090_n_spl_;
  wire g2091_n_spl_;
  wire g2092_n_spl_;
  wire g2092_n_spl_0;
  wire g2092_p_spl_;
  wire g2092_p_spl_0;
  wire g2094_n_spl_;
  wire g2094_p_spl_;
  wire g2095_n_spl_;
  wire g2095_p_spl_;
  wire g2089_n_spl_;
  wire g2097_p_spl_;
  wire g2089_p_spl_;
  wire g2097_n_spl_;
  wire g2098_n_spl_;
  wire g2098_p_spl_;
  wire g2088_n_spl_;
  wire g2100_p_spl_;
  wire g2088_p_spl_;
  wire g2100_n_spl_;
  wire g2101_n_spl_;
  wire g2101_p_spl_;
  wire g2087_n_spl_;
  wire g2103_p_spl_;
  wire g2087_p_spl_;
  wire g2103_n_spl_;
  wire g2104_n_spl_;
  wire g2104_p_spl_;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_01;
  wire G14_p_spl_1;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_1;
  wire g2112_p_spl_;
  wire g2113_p_spl_;
  wire g2112_n_spl_;
  wire g2113_n_spl_;
  wire g2114_n_spl_;
  wire g2114_n_spl_0;
  wire g2114_p_spl_;
  wire g2114_p_spl_0;
  wire g2116_n_spl_;
  wire g2116_p_spl_;
  wire g2117_n_spl_;
  wire g2117_p_spl_;
  wire g2111_n_spl_;
  wire g2119_p_spl_;
  wire g2111_p_spl_;
  wire g2119_n_spl_;
  wire g2120_n_spl_;
  wire g2120_p_spl_;
  wire g2110_n_spl_;
  wire g2122_p_spl_;
  wire g2110_p_spl_;
  wire g2122_n_spl_;
  wire g2123_n_spl_;
  wire g2123_p_spl_;
  wire g2109_n_spl_;
  wire g2125_p_spl_;
  wire g2109_p_spl_;
  wire g2125_n_spl_;
  wire g2126_n_spl_;
  wire g2126_p_spl_;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_1;
  wire g2134_p_spl_;
  wire g2135_p_spl_;
  wire g2134_n_spl_;
  wire g2135_n_spl_;
  wire g2136_n_spl_;
  wire g2136_n_spl_0;
  wire g2136_p_spl_;
  wire g2136_p_spl_0;
  wire g2138_n_spl_;
  wire g2138_p_spl_;
  wire g2139_n_spl_;
  wire g2139_p_spl_;
  wire g2133_n_spl_;
  wire g2141_p_spl_;
  wire g2133_p_spl_;
  wire g2141_n_spl_;
  wire g2142_n_spl_;
  wire g2142_p_spl_;
  wire g2132_n_spl_;
  wire g2144_p_spl_;
  wire g2132_p_spl_;
  wire g2144_n_spl_;
  wire g2145_n_spl_;
  wire g2145_p_spl_;
  wire g2131_n_spl_;
  wire g2147_p_spl_;
  wire g2131_p_spl_;
  wire g2147_n_spl_;
  wire g2148_n_spl_;
  wire g2148_p_spl_;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire g2156_p_spl_;
  wire g2157_p_spl_;
  wire g2156_n_spl_;
  wire g2157_n_spl_;
  wire g2158_n_spl_;
  wire g2158_p_spl_;
  wire g2160_n_spl_;
  wire g2160_p_spl_;
  wire g2161_n_spl_;
  wire g2161_p_spl_;
  wire g2155_n_spl_;
  wire g2163_p_spl_;
  wire g2155_p_spl_;
  wire g2163_n_spl_;
  wire g2164_n_spl_;
  wire g2164_p_spl_;
  wire g2154_n_spl_;
  wire g2166_p_spl_;
  wire g2154_p_spl_;
  wire g2166_n_spl_;
  wire g2167_n_spl_;
  wire g2167_p_spl_;
  wire g2153_n_spl_;
  wire g2169_p_spl_;
  wire g2153_p_spl_;
  wire g2169_n_spl_;
  wire g2170_n_spl_;
  wire g2170_p_spl_;
  wire g2177_p_spl_;
  wire g2177_n_spl_;
  wire g2178_p_spl_;
  wire g2179_n_spl_;
  wire g2178_n_spl_;
  wire g2179_p_spl_;
  wire g2180_n_spl_;
  wire g2180_p_spl_;
  wire g2176_n_spl_;
  wire g2182_p_spl_;
  wire g2176_p_spl_;
  wire g2182_n_spl_;
  wire g2183_n_spl_;
  wire g2183_p_spl_;
  wire g2175_n_spl_;
  wire g2185_p_spl_;
  wire g2175_p_spl_;
  wire g2185_n_spl_;
  wire g2186_n_spl_;
  wire g2186_p_spl_;
  wire g2192_n_spl_;
  wire g2193_n_spl_;
  wire g2192_p_spl_;
  wire g2193_p_spl_;
  wire g2194_n_spl_;
  wire g2191_n_spl_;
  wire g2196_p_spl_;
  wire g2191_p_spl_;
  wire g2196_n_spl_;
  wire g2197_n_spl_;
  wire g2201_n_spl_;
  wire g2203_p_spl_;
  wire g2201_p_spl_;
  wire g2203_n_spl_;
  wire g2204_n_spl_;
  wire g2204_p_spl_;
  wire g2205_n_spl_;
  wire g2207_p_spl_;
  wire g2208_n_spl_;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_000;
  wire G21_p_spl_001;
  wire G21_p_spl_01;
  wire G21_p_spl_010;
  wire G21_p_spl_011;
  wire G21_p_spl_1;
  wire G21_p_spl_10;
  wire G21_p_spl_100;
  wire G21_p_spl_101;
  wire G21_p_spl_11;
  wire g1631_p_spl_;
  wire g2228_n_spl_;
  wire g2230_p_spl_;
  wire g1975_n_spl_;
  wire g1997_n_spl_;
  wire g2019_n_spl_;
  wire g2041_n_spl_;
  wire g2063_n_spl_;
  wire g2085_n_spl_;
  wire g2107_n_spl_;
  wire g2129_n_spl_;
  wire g2151_n_spl_;
  wire g2173_n_spl_;
  wire g2189_n_spl_;
  wire g2200_n_spl_;
  wire g2212_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    n2491_lo_p,
    n2491_lo
  );


  not

  (
    n2491_lo_n,
    n2491_lo
  );


  buf

  (
    n2599_lo_p,
    n2599_lo
  );


  not

  (
    n2599_lo_n,
    n2599_lo
  );


  buf

  (
    n2611_lo_p,
    n2611_lo
  );


  not

  (
    n2611_lo_n,
    n2611_lo
  );


  buf

  (
    n2623_lo_p,
    n2623_lo
  );


  not

  (
    n2623_lo_n,
    n2623_lo
  );


  buf

  (
    n2635_lo_p,
    n2635_lo
  );


  not

  (
    n2635_lo_n,
    n2635_lo
  );


  buf

  (
    n2647_lo_p,
    n2647_lo
  );


  not

  (
    n2647_lo_n,
    n2647_lo
  );


  buf

  (
    n2659_lo_p,
    n2659_lo
  );


  not

  (
    n2659_lo_n,
    n2659_lo
  );


  buf

  (
    n2671_lo_p,
    n2671_lo
  );


  not

  (
    n2671_lo_n,
    n2671_lo
  );


  buf

  (
    n2683_lo_p,
    n2683_lo
  );


  not

  (
    n2683_lo_n,
    n2683_lo
  );


  buf

  (
    n2734_lo_p,
    n2734_lo
  );


  not

  (
    n2734_lo_n,
    n2734_lo
  );


  buf

  (
    n2746_lo_p,
    n2746_lo
  );


  not

  (
    n2746_lo_n,
    n2746_lo
  );


  buf

  (
    n2758_lo_p,
    n2758_lo
  );


  not

  (
    n2758_lo_n,
    n2758_lo
  );


  buf

  (
    n2770_lo_p,
    n2770_lo
  );


  not

  (
    n2770_lo_n,
    n2770_lo
  );


  buf

  (
    n2782_lo_p,
    n2782_lo
  );


  not

  (
    n2782_lo_n,
    n2782_lo
  );


  buf

  (
    n2794_lo_p,
    n2794_lo
  );


  not

  (
    n2794_lo_n,
    n2794_lo
  );


  buf

  (
    n2797_lo_p,
    n2797_lo
  );


  not

  (
    n2797_lo_n,
    n2797_lo
  );


  buf

  (
    n2806_lo_p,
    n2806_lo
  );


  not

  (
    n2806_lo_n,
    n2806_lo
  );


  buf

  (
    n2809_lo_p,
    n2809_lo
  );


  not

  (
    n2809_lo_n,
    n2809_lo
  );


  buf

  (
    n2818_lo_p,
    n2818_lo
  );


  not

  (
    n2818_lo_n,
    n2818_lo
  );


  buf

  (
    n2821_lo_p,
    n2821_lo
  );


  not

  (
    n2821_lo_n,
    n2821_lo
  );


  buf

  (
    n2830_lo_p,
    n2830_lo
  );


  not

  (
    n2830_lo_n,
    n2830_lo
  );


  buf

  (
    n2833_lo_p,
    n2833_lo
  );


  not

  (
    n2833_lo_n,
    n2833_lo
  );


  buf

  (
    n2839_lo_p,
    n2839_lo
  );


  not

  (
    n2839_lo_n,
    n2839_lo
  );


  buf

  (
    n2842_lo_p,
    n2842_lo
  );


  not

  (
    n2842_lo_n,
    n2842_lo
  );


  buf

  (
    n2845_lo_p,
    n2845_lo
  );


  not

  (
    n2845_lo_n,
    n2845_lo
  );


  buf

  (
    n2848_lo_p,
    n2848_lo
  );


  not

  (
    n2848_lo_n,
    n2848_lo
  );


  buf

  (
    n2851_lo_p,
    n2851_lo
  );


  not

  (
    n2851_lo_n,
    n2851_lo
  );


  buf

  (
    n2854_lo_p,
    n2854_lo
  );


  not

  (
    n2854_lo_n,
    n2854_lo
  );


  buf

  (
    n2857_lo_p,
    n2857_lo
  );


  not

  (
    n2857_lo_n,
    n2857_lo
  );


  buf

  (
    n2860_lo_p,
    n2860_lo
  );


  not

  (
    n2860_lo_n,
    n2860_lo
  );


  buf

  (
    n2863_lo_p,
    n2863_lo
  );


  not

  (
    n2863_lo_n,
    n2863_lo
  );


  buf

  (
    n3737_o2_p,
    n3737_o2
  );


  not

  (
    n3737_o2_n,
    n3737_o2
  );


  buf

  (
    n3736_o2_p,
    n3736_o2
  );


  not

  (
    n3736_o2_n,
    n3736_o2
  );


  buf

  (
    n3801_o2_p,
    n3801_o2
  );


  not

  (
    n3801_o2_n,
    n3801_o2
  );


  buf

  (
    n3836_o2_p,
    n3836_o2
  );


  not

  (
    n3836_o2_n,
    n3836_o2
  );


  buf

  (
    n3885_o2_p,
    n3885_o2
  );


  not

  (
    n3885_o2_n,
    n3885_o2
  );


  buf

  (
    n3902_o2_p,
    n3902_o2
  );


  not

  (
    n3902_o2_n,
    n3902_o2
  );


  buf

  (
    n4002_o2_p,
    n4002_o2
  );


  not

  (
    n4002_o2_n,
    n4002_o2
  );


  buf

  (
    n4052_o2_p,
    n4052_o2
  );


  not

  (
    n4052_o2_n,
    n4052_o2
  );


  buf

  (
    n4067_o2_p,
    n4067_o2
  );


  not

  (
    n4067_o2_n,
    n4067_o2
  );


  buf

  (
    n4162_o2_p,
    n4162_o2
  );


  not

  (
    n4162_o2_n,
    n4162_o2
  );


  buf

  (
    n4212_o2_p,
    n4212_o2
  );


  not

  (
    n4212_o2_n,
    n4212_o2
  );


  buf

  (
    n4227_o2_p,
    n4227_o2
  );


  not

  (
    n4227_o2_n,
    n4227_o2
  );


  buf

  (
    n4321_o2_p,
    n4321_o2
  );


  not

  (
    n4321_o2_n,
    n4321_o2
  );


  buf

  (
    n4367_o2_p,
    n4367_o2
  );


  not

  (
    n4367_o2_n,
    n4367_o2
  );


  buf

  (
    n4383_o2_p,
    n4383_o2
  );


  not

  (
    n4383_o2_n,
    n4383_o2
  );


  buf

  (
    n4475_o2_p,
    n4475_o2
  );


  not

  (
    n4475_o2_n,
    n4475_o2
  );


  buf

  (
    n4523_o2_p,
    n4523_o2
  );


  not

  (
    n4523_o2_n,
    n4523_o2
  );


  buf

  (
    n4537_o2_p,
    n4537_o2
  );


  not

  (
    n4537_o2_n,
    n4537_o2
  );


  buf

  (
    n4628_o2_p,
    n4628_o2
  );


  not

  (
    n4628_o2_n,
    n4628_o2
  );


  buf

  (
    n4674_o2_p,
    n4674_o2
  );


  not

  (
    n4674_o2_n,
    n4674_o2
  );


  buf

  (
    n4688_o2_p,
    n4688_o2
  );


  not

  (
    n4688_o2_n,
    n4688_o2
  );


  buf

  (
    n4791_o2_p,
    n4791_o2
  );


  not

  (
    n4791_o2_n,
    n4791_o2
  );


  buf

  (
    n4835_o2_p,
    n4835_o2
  );


  not

  (
    n4835_o2_n,
    n4835_o2
  );


  buf

  (
    n4868_o2_p,
    n4868_o2
  );


  not

  (
    n4868_o2_n,
    n4868_o2
  );


  buf

  (
    n5086_o2_p,
    n5086_o2
  );


  not

  (
    n5086_o2_n,
    n5086_o2
  );


  buf

  (
    n5130_o2_p,
    n5130_o2
  );


  not

  (
    n5130_o2_n,
    n5130_o2
  );


  buf

  (
    n5188_o2_p,
    n5188_o2
  );


  not

  (
    n5188_o2_n,
    n5188_o2
  );


  buf

  (
    n5402_o2_p,
    n5402_o2
  );


  not

  (
    n5402_o2_n,
    n5402_o2
  );


  buf

  (
    n5445_o2_p,
    n5445_o2
  );


  not

  (
    n5445_o2_n,
    n5445_o2
  );


  buf

  (
    n5500_o2_p,
    n5500_o2
  );


  not

  (
    n5500_o2_n,
    n5500_o2
  );


  buf

  (
    n5707_o2_p,
    n5707_o2
  );


  not

  (
    n5707_o2_n,
    n5707_o2
  );


  buf

  (
    n5745_o2_p,
    n5745_o2
  );


  not

  (
    n5745_o2_n,
    n5745_o2
  );


  buf

  (
    n5801_o2_p,
    n5801_o2
  );


  not

  (
    n5801_o2_n,
    n5801_o2
  );


  buf

  (
    n4836_o2_p,
    n4836_o2
  );


  not

  (
    n4836_o2_n,
    n4836_o2
  );


  buf

  (
    n4837_o2_p,
    n4837_o2
  );


  not

  (
    n4837_o2_n,
    n4837_o2
  );


  buf

  (
    n4838_o2_p,
    n4838_o2
  );


  not

  (
    n4838_o2_n,
    n4838_o2
  );


  buf

  (
    n4839_o2_p,
    n4839_o2
  );


  not

  (
    n4839_o2_n,
    n4839_o2
  );


  buf

  (
    n4840_o2_p,
    n4840_o2
  );


  not

  (
    n4840_o2_n,
    n4840_o2
  );


  buf

  (
    n4841_o2_p,
    n4841_o2
  );


  not

  (
    n4841_o2_n,
    n4841_o2
  );


  buf

  (
    n4842_o2_p,
    n4842_o2
  );


  not

  (
    n4842_o2_n,
    n4842_o2
  );


  buf

  (
    n4843_o2_p,
    n4843_o2
  );


  not

  (
    n4843_o2_n,
    n4843_o2
  );


  buf

  (
    n4844_o2_p,
    n4844_o2
  );


  not

  (
    n4844_o2_n,
    n4844_o2
  );


  buf

  (
    n4845_o2_p,
    n4845_o2
  );


  not

  (
    n4845_o2_n,
    n4845_o2
  );


  buf

  (
    n4846_o2_p,
    n4846_o2
  );


  not

  (
    n4846_o2_n,
    n4846_o2
  );


  buf

  (
    n4847_o2_p,
    n4847_o2
  );


  not

  (
    n4847_o2_n,
    n4847_o2
  );


  buf

  (
    n4848_o2_p,
    n4848_o2
  );


  not

  (
    n4848_o2_n,
    n4848_o2
  );


  buf

  (
    n4849_o2_p,
    n4849_o2
  );


  not

  (
    n4849_o2_n,
    n4849_o2
  );


  buf

  (
    n4850_o2_p,
    n4850_o2
  );


  not

  (
    n4850_o2_n,
    n4850_o2
  );


  buf

  (
    n4867_o2_p,
    n4867_o2
  );


  not

  (
    n4867_o2_n,
    n4867_o2
  );


  buf

  (
    n4908_o2_p,
    n4908_o2
  );


  not

  (
    n4908_o2_n,
    n4908_o2
  );


  buf

  (
    n6081_o2_p,
    n6081_o2
  );


  not

  (
    n6081_o2_n,
    n6081_o2
  );


  buf

  (
    n6120_o2_p,
    n6120_o2
  );


  not

  (
    n6120_o2_n,
    n6120_o2
  );


  buf

  (
    n316_inv_p,
    n316_inv
  );


  not

  (
    n316_inv_n,
    n316_inv
  );


  buf

  (
    n4960_o2_p,
    n4960_o2
  );


  not

  (
    n4960_o2_n,
    n4960_o2
  );


  buf

  (
    n6203_o2_p,
    n6203_o2
  );


  not

  (
    n6203_o2_n,
    n6203_o2
  );


  buf

  (
    n325_inv_p,
    n325_inv
  );


  not

  (
    n325_inv_n,
    n325_inv
  );


  buf

  (
    n328_inv_p,
    n328_inv
  );


  not

  (
    n328_inv_n,
    n328_inv
  );


  buf

  (
    n331_inv_p,
    n331_inv
  );


  not

  (
    n331_inv_n,
    n331_inv
  );


  buf

  (
    n5189_o2_p,
    n5189_o2
  );


  not

  (
    n5189_o2_n,
    n5189_o2
  );


  buf

  (
    n6594_o2_p,
    n6594_o2
  );


  not

  (
    n6594_o2_n,
    n6594_o2
  );


  buf

  (
    n340_inv_p,
    n340_inv
  );


  not

  (
    n340_inv_n,
    n340_inv
  );


  buf

  (
    n6631_o2_p,
    n6631_o2
  );


  not

  (
    n6631_o2_n,
    n6631_o2
  );


  buf

  (
    n346_inv_p,
    n346_inv
  );


  not

  (
    n346_inv_n,
    n346_inv
  );


  buf

  (
    n5388_o2_p,
    n5388_o2
  );


  not

  (
    n5388_o2_n,
    n5388_o2
  );


  buf

  (
    n6725_o2_p,
    n6725_o2
  );


  not

  (
    n6725_o2_n,
    n6725_o2
  );


  buf

  (
    n355_inv_p,
    n355_inv
  );


  not

  (
    n355_inv_n,
    n355_inv
  );


  buf

  (
    n358_inv_p,
    n358_inv
  );


  not

  (
    n358_inv_n,
    n358_inv
  );


  buf

  (
    n5612_o2_p,
    n5612_o2
  );


  not

  (
    n5612_o2_n,
    n5612_o2
  );


  buf

  (
    n1127_o2_p,
    n1127_o2
  );


  not

  (
    n1127_o2_n,
    n1127_o2
  );


  buf

  (
    n367_inv_p,
    n367_inv
  );


  not

  (
    n367_inv_n,
    n367_inv
  );


  buf

  (
    n1231_o2_p,
    n1231_o2
  );


  not

  (
    n1231_o2_n,
    n1231_o2
  );


  buf

  (
    n373_inv_p,
    n373_inv
  );


  not

  (
    n373_inv_n,
    n373_inv
  );


  buf

  (
    n5802_o2_p,
    n5802_o2
  );


  not

  (
    n5802_o2_n,
    n5802_o2
  );


  buf

  (
    n1232_o2_p,
    n1232_o2
  );


  not

  (
    n1232_o2_n,
    n1232_o2
  );


  buf

  (
    n382_inv_p,
    n382_inv
  );


  not

  (
    n382_inv_n,
    n382_inv
  );


  buf

  (
    n385_inv_p,
    n385_inv
  );


  not

  (
    n385_inv_n,
    n385_inv
  );


  buf

  (
    n6023_o2_p,
    n6023_o2
  );


  not

  (
    n6023_o2_n,
    n6023_o2
  );


  buf

  (
    n1235_o2_p,
    n1235_o2
  );


  not

  (
    n1235_o2_n,
    n1235_o2
  );


  buf

  (
    n394_inv_p,
    n394_inv
  );


  not

  (
    n394_inv_n,
    n394_inv
  );


  buf

  (
    n1347_o2_p,
    n1347_o2
  );


  not

  (
    n1347_o2_n,
    n1347_o2
  );


  buf

  (
    n400_inv_p,
    n400_inv
  );


  not

  (
    n400_inv_n,
    n400_inv
  );


  buf

  (
    n6383_o2_p,
    n6383_o2
  );


  not

  (
    n6383_o2_n,
    n6383_o2
  );


  buf

  (
    n1348_o2_p,
    n1348_o2
  );


  not

  (
    n1348_o2_n,
    n1348_o2
  );


  buf

  (
    n409_inv_p,
    n409_inv
  );


  not

  (
    n409_inv_n,
    n409_inv
  );


  buf

  (
    n1351_o2_p,
    n1351_o2
  );


  not

  (
    n1351_o2_n,
    n1351_o2
  );


  buf

  (
    n1461_o2_p,
    n1461_o2
  );


  not

  (
    n1461_o2_n,
    n1461_o2
  );


  buf

  (
    n418_inv_p,
    n418_inv
  );


  not

  (
    n418_inv_n,
    n418_inv
  );


  buf

  (
    n6024_o2_p,
    n6024_o2
  );


  not

  (
    n6024_o2_n,
    n6024_o2
  );


  buf

  (
    n6025_o2_p,
    n6025_o2
  );


  not

  (
    n6025_o2_n,
    n6025_o2
  );


  buf

  (
    n6026_o2_p,
    n6026_o2
  );


  not

  (
    n6026_o2_n,
    n6026_o2
  );


  buf

  (
    n6027_o2_p,
    n6027_o2
  );


  not

  (
    n6027_o2_n,
    n6027_o2
  );


  buf

  (
    n6028_o2_p,
    n6028_o2
  );


  not

  (
    n6028_o2_n,
    n6028_o2
  );


  buf

  (
    n6029_o2_p,
    n6029_o2
  );


  not

  (
    n6029_o2_n,
    n6029_o2
  );


  buf

  (
    n6030_o2_p,
    n6030_o2
  );


  not

  (
    n6030_o2_n,
    n6030_o2
  );


  buf

  (
    n6031_o2_p,
    n6031_o2
  );


  not

  (
    n6031_o2_n,
    n6031_o2
  );


  buf

  (
    n6032_o2_p,
    n6032_o2
  );


  not

  (
    n6032_o2_n,
    n6032_o2
  );


  buf

  (
    n6033_o2_p,
    n6033_o2
  );


  not

  (
    n6033_o2_n,
    n6033_o2
  );


  buf

  (
    n6034_o2_p,
    n6034_o2
  );


  not

  (
    n6034_o2_n,
    n6034_o2
  );


  buf

  (
    n6035_o2_p,
    n6035_o2
  );


  not

  (
    n6035_o2_n,
    n6035_o2
  );


  buf

  (
    n6036_o2_p,
    n6036_o2
  );


  not

  (
    n6036_o2_n,
    n6036_o2
  );


  buf

  (
    n6037_o2_p,
    n6037_o2
  );


  not

  (
    n6037_o2_n,
    n6037_o2
  );


  buf

  (
    n6038_o2_p,
    n6038_o2
  );


  not

  (
    n6038_o2_n,
    n6038_o2
  );


  buf

  (
    n6053_o2_p,
    n6053_o2
  );


  not

  (
    n6053_o2_n,
    n6053_o2
  );


  buf

  (
    n6726_o2_p,
    n6726_o2
  );


  not

  (
    n6726_o2_n,
    n6726_o2
  );


  buf

  (
    n6148_o2_p,
    n6148_o2
  );


  not

  (
    n6148_o2_n,
    n6148_o2
  );


  buf

  (
    n1463_o2_p,
    n1463_o2
  );


  not

  (
    n1463_o2_n,
    n1463_o2
  );


  buf

  (
    n1573_o2_p,
    n1573_o2
  );


  not

  (
    n1573_o2_n,
    n1573_o2
  );


  buf

  (
    n481_inv_p,
    n481_inv
  );


  not

  (
    n481_inv_n,
    n481_inv
  );


  buf

  (
    n6201_o2_p,
    n6201_o2
  );


  not

  (
    n6201_o2_n,
    n6201_o2
  );


  buf

  (
    n487_inv_p,
    n487_inv
  );


  not

  (
    n487_inv_n,
    n487_inv
  );


  buf

  (
    n490_inv_p,
    n490_inv
  );


  not

  (
    n490_inv_n,
    n490_inv
  );


  buf

  (
    n493_inv_p,
    n493_inv
  );


  not

  (
    n493_inv_n,
    n493_inv
  );


  buf

  (
    n1574_o2_p,
    n1574_o2
  );


  not

  (
    n1574_o2_n,
    n1574_o2
  );


  buf

  (
    n499_inv_p,
    n499_inv
  );


  not

  (
    n499_inv_n,
    n499_inv
  );


  buf

  (
    n502_inv_p,
    n502_inv
  );


  not

  (
    n502_inv_n,
    n502_inv
  );


  buf

  (
    n772_o2_p,
    n772_o2
  );


  not

  (
    n772_o2_n,
    n772_o2
  );


  buf

  (
    n6482_o2_p,
    n6482_o2
  );


  not

  (
    n6482_o2_n,
    n6482_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    n1577_o2_p,
    n1577_o2
  );


  not

  (
    n1577_o2_n,
    n1577_o2
  );


  buf

  (
    n1678_o2_p,
    n1678_o2
  );


  not

  (
    n1678_o2_n,
    n1678_o2
  );


  buf

  (
    n520_inv_p,
    n520_inv
  );


  not

  (
    n520_inv_n,
    n520_inv
  );


  buf

  (
    n523_inv_p,
    n523_inv
  );


  not

  (
    n523_inv_n,
    n523_inv
  );


  buf

  (
    n6727_o2_p,
    n6727_o2
  );


  not

  (
    n6727_o2_n,
    n6727_o2
  );


  buf

  (
    n529_inv_p,
    n529_inv
  );


  not

  (
    n529_inv_n,
    n529_inv
  );


  buf

  (
    n1679_o2_p,
    n1679_o2
  );


  not

  (
    n1679_o2_n,
    n1679_o2
  );


  buf

  (
    n535_inv_p,
    n535_inv
  );


  not

  (
    n535_inv_n,
    n535_inv
  );


  buf

  (
    n848_o2_p,
    n848_o2
  );


  not

  (
    n848_o2_n,
    n848_o2
  );


  buf

  (
    n541_inv_p,
    n541_inv
  );


  not

  (
    n541_inv_n,
    n541_inv
  );


  buf

  (
    n544_inv_p,
    n544_inv
  );


  not

  (
    n544_inv_n,
    n544_inv
  );


  buf

  (
    lo110_buf_o2_p,
    lo110_buf_o2
  );


  not

  (
    lo110_buf_o2_n,
    lo110_buf_o2
  );


  buf

  (
    n1682_o2_p,
    n1682_o2
  );


  not

  (
    n1682_o2_n,
    n1682_o2
  );


  buf

  (
    n1775_o2_p,
    n1775_o2
  );


  not

  (
    n1775_o2_n,
    n1775_o2
  );


  buf

  (
    n512_o2_p,
    n512_o2
  );


  not

  (
    n512_o2_n,
    n512_o2
  );


  buf

  (
    n559_inv_p,
    n559_inv
  );


  not

  (
    n559_inv_n,
    n559_inv
  );


  buf

  (
    n562_inv_p,
    n562_inv
  );


  not

  (
    n562_inv_n,
    n562_inv
  );


  buf

  (
    n2210_o2_p,
    n2210_o2
  );


  not

  (
    n2210_o2_n,
    n2210_o2
  );


  buf

  (
    n2126_o2_p,
    n2126_o2
  );


  not

  (
    n2126_o2_n,
    n2126_o2
  );


  buf

  (
    n2010_o2_p,
    n2010_o2
  );


  not

  (
    n2010_o2_n,
    n2010_o2
  );


  buf

  (
    n1776_o2_p,
    n1776_o2
  );


  not

  (
    n1776_o2_n,
    n1776_o2
  );


  buf

  (
    n577_inv_p,
    n577_inv
  );


  not

  (
    n577_inv_n,
    n577_inv
  );


  buf

  (
    n580_inv_p,
    n580_inv
  );


  not

  (
    n580_inv_n,
    n580_inv
  );


  buf

  (
    n932_o2_p,
    n932_o2
  );


  not

  (
    n932_o2_n,
    n932_o2
  );


  buf

  (
    n548_o2_p,
    n548_o2
  );


  not

  (
    n548_o2_n,
    n548_o2
  );


  buf

  (
    lo114_buf_o2_p,
    lo114_buf_o2
  );


  not

  (
    lo114_buf_o2_n,
    lo114_buf_o2
  );


  buf

  (
    n1779_o2_p,
    n1779_o2
  );


  not

  (
    n1779_o2_n,
    n1779_o2
  );


  buf

  (
    n1864_o2_p,
    n1864_o2
  );


  not

  (
    n1864_o2_n,
    n1864_o2
  );


  buf

  (
    n598_inv_p,
    n598_inv
  );


  not

  (
    n598_inv_n,
    n598_inv
  );


  buf

  (
    n601_inv_p,
    n601_inv
  );


  not

  (
    n601_inv_n,
    n601_inv
  );


  buf

  (
    n592_o2_p,
    n592_o2
  );


  not

  (
    n592_o2_n,
    n592_o2
  );


  buf

  (
    lo010_buf_o2_p,
    lo010_buf_o2
  );


  not

  (
    lo010_buf_o2_n,
    lo010_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo018_buf_o2_p,
    lo018_buf_o2
  );


  not

  (
    lo018_buf_o2_n,
    lo018_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo026_buf_o2_p,
    lo026_buf_o2
  );


  not

  (
    lo026_buf_o2_n,
    lo026_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo034_buf_o2_p,
    lo034_buf_o2
  );


  not

  (
    lo034_buf_o2_n,
    lo034_buf_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo046_buf_o2_p,
    lo046_buf_o2
  );


  not

  (
    lo046_buf_o2_n,
    lo046_buf_o2
  );


  buf

  (
    lo050_buf_o2_p,
    lo050_buf_o2
  );


  not

  (
    lo050_buf_o2_n,
    lo050_buf_o2
  );


  buf

  (
    lo054_buf_o2_p,
    lo054_buf_o2
  );


  not

  (
    lo054_buf_o2_n,
    lo054_buf_o2
  );


  buf

  (
    lo058_buf_o2_p,
    lo058_buf_o2
  );


  not

  (
    lo058_buf_o2_n,
    lo058_buf_o2
  );


  buf

  (
    lo062_buf_o2_p,
    lo062_buf_o2
  );


  not

  (
    lo062_buf_o2_n,
    lo062_buf_o2
  );


  buf

  (
    lo066_buf_o2_p,
    lo066_buf_o2
  );


  not

  (
    lo066_buf_o2_n,
    lo066_buf_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    n655_inv_p,
    n655_inv
  );


  not

  (
    n655_inv_n,
    n655_inv
  );


  buf

  (
    n2013_o2_p,
    n2013_o2
  );


  not

  (
    n2013_o2_n,
    n2013_o2
  );


  buf

  (
    n2129_o2_p,
    n2129_o2
  );


  not

  (
    n2129_o2_n,
    n2129_o2
  );


  buf

  (
    n2213_o2_p,
    n2213_o2
  );


  not

  (
    n2213_o2_n,
    n2213_o2
  );


  buf

  (
    n2243_o2_p,
    n2243_o2
  );


  not

  (
    n2243_o2_n,
    n2243_o2
  );


  buf

  (
    n2175_o2_p,
    n2175_o2
  );


  not

  (
    n2175_o2_n,
    n2175_o2
  );


  buf

  (
    n2075_o2_p,
    n2075_o2
  );


  not

  (
    n2075_o2_n,
    n2075_o2
  );


  buf

  (
    n1943_o2_p,
    n1943_o2
  );


  not

  (
    n1943_o2_n,
    n1943_o2
  );


  buf

  (
    n1865_o2_p,
    n1865_o2
  );


  not

  (
    n1865_o2_n,
    n1865_o2
  );


  buf

  (
    n682_inv_p,
    n682_inv
  );


  not

  (
    n682_inv_n,
    n682_inv
  );


  buf

  (
    lo094_buf_o2_p,
    lo094_buf_o2
  );


  not

  (
    lo094_buf_o2_n,
    lo094_buf_o2
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    n691_inv_p,
    n691_inv
  );


  not

  (
    n691_inv_n,
    n691_inv
  );


  buf

  (
    n451_o2_p,
    n451_o2
  );


  not

  (
    n451_o2_n,
    n451_o2
  );


  buf

  (
    n1024_o2_p,
    n1024_o2
  );


  not

  (
    n1024_o2_n,
    n1024_o2
  );


  buf

  (
    n700_inv_p,
    n700_inv
  );


  not

  (
    n700_inv_n,
    n700_inv
  );


  buf

  (
    n703_inv_p,
    n703_inv
  );


  not

  (
    n703_inv_n,
    n703_inv
  );


  buf

  (
    n706_inv_p,
    n706_inv
  );


  not

  (
    n706_inv_n,
    n706_inv
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    n1868_o2_p,
    n1868_o2
  );


  not

  (
    n1868_o2_n,
    n1868_o2
  );


  buf

  (
    n1945_o2_p,
    n1945_o2
  );


  not

  (
    n1945_o2_n,
    n1945_o2
  );


  buf

  (
    n718_inv_p,
    n718_inv
  );


  not

  (
    n718_inv_n,
    n718_inv
  );


  buf

  (
    n2045_o2_p,
    n2045_o2
  );


  not

  (
    n2045_o2_n,
    n2045_o2
  );


  buf

  (
    n1913_o2_p,
    n1913_o2
  );


  not

  (
    n1913_o2_n,
    n1913_o2
  );


  buf

  (
    n1749_o2_p,
    n1749_o2
  );


  not

  (
    n1749_o2_n,
    n1749_o2
  );


  buf

  (
    n1553_o2_p,
    n1553_o2
  );


  not

  (
    n1553_o2_n,
    n1553_o2
  );


  buf

  (
    n644_o2_p,
    n644_o2
  );


  not

  (
    n644_o2_n,
    n644_o2
  );


  buf

  (
    n736_inv_p,
    n736_inv
  );


  not

  (
    n736_inv_n,
    n736_inv
  );


  buf

  (
    lo098_buf_o2_p,
    lo098_buf_o2
  );


  not

  (
    lo098_buf_o2_n,
    lo098_buf_o2
  );


  buf

  (
    n1121_o2_p,
    n1121_o2
  );


  not

  (
    n1121_o2_n,
    n1121_o2
  );


  buf

  (
    n1719_o2_p,
    n1719_o2
  );


  not

  (
    n1719_o2_n,
    n1719_o2
  );


  buf

  (
    n1523_o2_p,
    n1523_o2
  );


  not

  (
    n1523_o2_n,
    n1523_o2
  );


  buf

  (
    n464_o2_p,
    n464_o2
  );


  not

  (
    n464_o2_n,
    n464_o2
  );


  buf

  (
    n754_inv_p,
    n754_inv
  );


  not

  (
    n754_inv_n,
    n754_inv
  );


  buf

  (
    n757_inv_p,
    n757_inv
  );


  not

  (
    n757_inv_n,
    n757_inv
  );


  buf

  (
    n760_inv_p,
    n760_inv
  );


  not

  (
    n760_inv_n,
    n760_inv
  );


  buf

  (
    n2078_o2_p,
    n2078_o2
  );


  not

  (
    n2078_o2_n,
    n2078_o2
  );


  buf

  (
    n2079_o2_p,
    n2079_o2
  );


  not

  (
    n2079_o2_n,
    n2079_o2
  );


  buf

  (
    n2178_o2_p,
    n2178_o2
  );


  not

  (
    n2178_o2_n,
    n2178_o2
  );


  buf

  (
    n2179_o2_p,
    n2179_o2
  );


  not

  (
    n2179_o2_n,
    n2179_o2
  );


  buf

  (
    n2246_o2_p,
    n2246_o2
  );


  not

  (
    n2246_o2_n,
    n2246_o2
  );


  buf

  (
    n2247_o2_p,
    n2247_o2
  );


  not

  (
    n2247_o2_n,
    n2247_o2
  );


  buf

  (
    n2216_o2_p,
    n2216_o2
  );


  not

  (
    n2216_o2_n,
    n2216_o2
  );


  buf

  (
    n2217_o2_p,
    n2217_o2
  );


  not

  (
    n2217_o2_n,
    n2217_o2
  );


  buf

  (
    n2132_o2_p,
    n2132_o2
  );


  not

  (
    n2132_o2_n,
    n2132_o2
  );


  buf

  (
    n2133_o2_p,
    n2133_o2
  );


  not

  (
    n2133_o2_n,
    n2133_o2
  );


  buf

  (
    n2016_o2_p,
    n2016_o2
  );


  not

  (
    n2016_o2_n,
    n2016_o2
  );


  buf

  (
    n2017_o2_p,
    n2017_o2
  );


  not

  (
    n2017_o2_n,
    n2017_o2
  );


  buf

  (
    n1946_o2_p,
    n1946_o2
  );


  not

  (
    n1946_o2_n,
    n1946_o2
  );


  buf

  (
    n1556_o2_p,
    n1556_o2
  );


  not

  (
    n1556_o2_n,
    n1556_o2
  );


  buf

  (
    n1752_o2_p,
    n1752_o2
  );


  not

  (
    n1752_o2_n,
    n1752_o2
  );


  buf

  (
    n1916_o2_p,
    n1916_o2
  );


  not

  (
    n1916_o2_n,
    n1916_o2
  );


  buf

  (
    n2048_o2_p,
    n2048_o2
  );


  not

  (
    n2048_o2_n,
    n2048_o2
  );


  buf

  (
    n2102_o2_p,
    n2102_o2
  );


  not

  (
    n2102_o2_n,
    n2102_o2
  );


  buf

  (
    n1226_o2_p,
    n1226_o2
  );


  not

  (
    n1226_o2_n,
    n1226_o2
  );


  buf

  (
    n1986_o2_p,
    n1986_o2
  );


  not

  (
    n1986_o2_n,
    n1986_o2
  );


  buf

  (
    n1838_o2_p,
    n1838_o2
  );


  not

  (
    n1838_o2_n,
    n1838_o2
  );


  buf

  (
    n1658_o2_p,
    n1658_o2
  );


  not

  (
    n1658_o2_n,
    n1658_o2
  );


  buf

  (
    n829_inv_p,
    n829_inv
  );


  not

  (
    n829_inv_n,
    n829_inv
  );


  buf

  (
    n1526_o2_p,
    n1526_o2
  );


  not

  (
    n1526_o2_n,
    n1526_o2
  );


  buf

  (
    n1722_o2_p,
    n1722_o2
  );


  not

  (
    n1722_o2_n,
    n1722_o2
  );


  buf

  (
    n1808_o2_p,
    n1808_o2
  );


  not

  (
    n1808_o2_n,
    n1808_o2
  );


  buf

  (
    n1628_o2_p,
    n1628_o2
  );


  not

  (
    n1628_o2_n,
    n1628_o2
  );


  buf

  (
    n844_inv_p,
    n844_inv
  );


  not

  (
    n844_inv_n,
    n844_inv
  );


  buf

  (
    n847_inv_p,
    n847_inv
  );


  not

  (
    n847_inv_n,
    n847_inv
  );


  buf

  (
    n1583_o2_p,
    n1583_o2
  );


  not

  (
    n1583_o2_n,
    n1583_o2
  );


  buf

  (
    n1787_o2_p,
    n1787_o2
  );


  not

  (
    n1787_o2_n,
    n1787_o2
  );


  buf

  (
    n1959_o2_p,
    n1959_o2
  );


  not

  (
    n1959_o2_n,
    n1959_o2
  );


  buf

  (
    n2099_o2_p,
    n2099_o2
  );


  not

  (
    n2099_o2_n,
    n2099_o2
  );


  buf

  (
    n2033_o2_p,
    n2033_o2
  );


  not

  (
    n2033_o2_n,
    n2033_o2
  );


  buf

  (
    n1877_o2_p,
    n1877_o2
  );


  not

  (
    n1877_o2_n,
    n1877_o2
  );


  buf

  (
    n1689_o2_p,
    n1689_o2
  );


  not

  (
    n1689_o2_n,
    n1689_o2
  );


  buf

  (
    n1355_o2_p,
    n1355_o2
  );


  not

  (
    n1355_o2_n,
    n1355_o2
  );


  buf

  (
    n1469_o2_p,
    n1469_o2
  );


  not

  (
    n1469_o2_n,
    n1469_o2
  );


  buf

  (
    n1238_o2_p,
    n1238_o2
  );


  not

  (
    n1238_o2_n,
    n1238_o2
  );


  buf

  (
    n1227_o2_p,
    n1227_o2
  );


  not

  (
    n1227_o2_n,
    n1227_o2
  );


  buf

  (
    n1124_o2_p,
    n1124_o2
  );


  not

  (
    n1124_o2_n,
    n1124_o2
  );


  buf

  (
    n704_o2_p,
    n704_o2
  );


  not

  (
    n704_o2_n,
    n704_o2
  );


  buf

  (
    n484_o2_p,
    n484_o2
  );


  not

  (
    n484_o2_n,
    n484_o2
  );


  buf

  (
    n1338_o2_p,
    n1338_o2
  );


  not

  (
    n1338_o2_n,
    n1338_o2
  );


  buf

  (
    n1449_o2_p,
    n1449_o2
  );


  not

  (
    n1449_o2_n,
    n1449_o2
  );


  buf

  (
    n1558_o2_p,
    n1558_o2
  );


  not

  (
    n1558_o2_n,
    n1558_o2
  );


  buf

  (
    n1754_o2_p,
    n1754_o2
  );


  not

  (
    n1754_o2_n,
    n1754_o2
  );


  buf

  (
    n1918_o2_p,
    n1918_o2
  );


  not

  (
    n1918_o2_n,
    n1918_o2
  );


  buf

  (
    n2050_o2_p,
    n2050_o2
  );


  not

  (
    n2050_o2_n,
    n2050_o2
  );


  buf

  (
    n2104_o2_p,
    n2104_o2
  );


  not

  (
    n2104_o2_n,
    n2104_o2
  );


  buf

  (
    n1988_o2_p,
    n1988_o2
  );


  not

  (
    n1988_o2_n,
    n1988_o2
  );


  buf

  (
    n1840_o2_p,
    n1840_o2
  );


  not

  (
    n1840_o2_n,
    n1840_o2
  );


  buf

  (
    n1660_o2_p,
    n1660_o2
  );


  not

  (
    n1660_o2_n,
    n1660_o2
  );


  buf

  (
    n708_o2_p,
    n708_o2
  );


  not

  (
    n708_o2_n,
    n708_o2
  );


  buf

  (
    n768_o2_p,
    n768_o2
  );


  not

  (
    n768_o2_n,
    n768_o2
  );


  buf

  (
    lo102_buf_o2_p,
    lo102_buf_o2
  );


  not

  (
    lo102_buf_o2_n,
    lo102_buf_o2
  );


  buf

  (
    n1631_o2_p,
    n1631_o2
  );


  not

  (
    n1631_o2_n,
    n1631_o2
  );


  buf

  (
    n1632_o2_p,
    n1632_o2
  );


  not

  (
    n1632_o2_n,
    n1632_o2
  );


  buf

  (
    n1811_o2_p,
    n1811_o2
  );


  not

  (
    n1811_o2_n,
    n1811_o2
  );


  buf

  (
    n1812_o2_p,
    n1812_o2
  );


  not

  (
    n1812_o2_n,
    n1812_o2
  );


  buf

  (
    n1889_o2_p,
    n1889_o2
  );


  not

  (
    n1889_o2_n,
    n1889_o2
  );


  buf

  (
    n1890_o2_p,
    n1890_o2
  );


  not

  (
    n1890_o2_n,
    n1890_o2
  );


  buf

  (
    n1725_o2_p,
    n1725_o2
  );


  not

  (
    n1725_o2_n,
    n1725_o2
  );


  buf

  (
    n1726_o2_p,
    n1726_o2
  );


  not

  (
    n1726_o2_n,
    n1726_o2
  );


  buf

  (
    n917_o2_p,
    n917_o2
  );


  not

  (
    n917_o2_n,
    n917_o2
  );


  buf

  (
    n918_o2_p,
    n918_o2
  );


  not

  (
    n918_o2_n,
    n918_o2
  );


  buf

  (
    n1003_o2_p,
    n1003_o2
  );


  not

  (
    n1003_o2_n,
    n1003_o2
  );


  buf

  (
    n1004_o2_p,
    n1004_o2
  );


  not

  (
    n1004_o2_n,
    n1004_o2
  );


  buf

  (
    n1097_o2_p,
    n1097_o2
  );


  not

  (
    n1097_o2_n,
    n1097_o2
  );


  buf

  (
    n1098_o2_p,
    n1098_o2
  );


  not

  (
    n1098_o2_n,
    n1098_o2
  );


  buf

  (
    n1199_o2_p,
    n1199_o2
  );


  not

  (
    n1199_o2_n,
    n1199_o2
  );


  buf

  (
    n1200_o2_p,
    n1200_o2
  );


  not

  (
    n1200_o2_n,
    n1200_o2
  );


  buf

  (
    n1309_o2_p,
    n1309_o2
  );


  not

  (
    n1309_o2_n,
    n1309_o2
  );


  buf

  (
    n1310_o2_p,
    n1310_o2
  );


  not

  (
    n1310_o2_n,
    n1310_o2
  );


  buf

  (
    n1420_o2_p,
    n1420_o2
  );


  not

  (
    n1420_o2_n,
    n1420_o2
  );


  buf

  (
    n1421_o2_p,
    n1421_o2
  );


  not

  (
    n1421_o2_n,
    n1421_o2
  );


  buf

  (
    n1529_o2_p,
    n1529_o2
  );


  not

  (
    n1529_o2_n,
    n1529_o2
  );


  buf

  (
    n1530_o2_p,
    n1530_o2
  );


  not

  (
    n1530_o2_n,
    n1530_o2
  );


  buf

  (
    n839_o2_p,
    n839_o2
  );


  not

  (
    n839_o2_n,
    n839_o2
  );


  buf

  (
    n840_o2_p,
    n840_o2
  );


  not

  (
    n840_o2_n,
    n840_o2
  );


  buf

  (
    n577_o2_p,
    n577_o2
  );


  not

  (
    n577_o2_n,
    n577_o2
  );


  buf

  (
    n623_o2_p,
    n623_o2
  );


  not

  (
    n623_o2_n,
    n623_o2
  );


  buf

  (
    n677_o2_p,
    n677_o2
  );


  not

  (
    n677_o2_n,
    n677_o2
  );


  buf

  (
    n739_o2_p,
    n739_o2
  );


  not

  (
    n739_o2_n,
    n739_o2
  );


  buf

  (
    n809_o2_p,
    n809_o2
  );


  not

  (
    n809_o2_n,
    n809_o2
  );


  buf

  (
    n887_o2_p,
    n887_o2
  );


  not

  (
    n887_o2_n,
    n887_o2
  );


  buf

  (
    n973_o2_p,
    n973_o2
  );


  not

  (
    n973_o2_n,
    n973_o2
  );


  buf

  (
    n1067_o2_p,
    n1067_o2
  );


  not

  (
    n1067_o2_n,
    n1067_o2
  );


  buf

  (
    n1169_o2_p,
    n1169_o2
  );


  not

  (
    n1169_o2_n,
    n1169_o2
  );


  buf

  (
    n1279_o2_p,
    n1279_o2
  );


  not

  (
    n1279_o2_n,
    n1279_o2
  );


  buf

  (
    n1390_o2_p,
    n1390_o2
  );


  not

  (
    n1390_o2_n,
    n1390_o2
  );


  buf

  (
    n1499_o2_p,
    n1499_o2
  );


  not

  (
    n1499_o2_n,
    n1499_o2
  );


  buf

  (
    n539_o2_p,
    n539_o2
  );


  not

  (
    n539_o2_n,
    n539_o2
  );


  buf

  (
    lo082_buf_o2_p,
    lo082_buf_o2
  );


  not

  (
    lo082_buf_o2_n,
    lo082_buf_o2
  );


  buf

  (
    n555_o2_p,
    n555_o2
  );


  not

  (
    n555_o2_n,
    n555_o2
  );


  buf

  (
    n601_o2_p,
    n601_o2
  );


  not

  (
    n601_o2_n,
    n601_o2
  );


  buf

  (
    n655_o2_p,
    n655_o2
  );


  not

  (
    n655_o2_n,
    n655_o2
  );


  buf

  (
    n717_o2_p,
    n717_o2
  );


  not

  (
    n717_o2_n,
    n717_o2
  );


  buf

  (
    n787_o2_p,
    n787_o2
  );


  not

  (
    n787_o2_n,
    n787_o2
  );


  buf

  (
    n865_o2_p,
    n865_o2
  );


  not

  (
    n865_o2_n,
    n865_o2
  );


  buf

  (
    n951_o2_p,
    n951_o2
  );


  not

  (
    n951_o2_n,
    n951_o2
  );


  buf

  (
    n1045_o2_p,
    n1045_o2
  );


  not

  (
    n1045_o2_n,
    n1045_o2
  );


  buf

  (
    n1147_o2_p,
    n1147_o2
  );


  not

  (
    n1147_o2_n,
    n1147_o2
  );


  buf

  (
    n1257_o2_p,
    n1257_o2
  );


  not

  (
    n1257_o2_n,
    n1257_o2
  );


  buf

  (
    n1374_o2_p,
    n1374_o2
  );


  not

  (
    n1374_o2_n,
    n1374_o2
  );


  buf

  (
    n1488_o2_p,
    n1488_o2
  );


  not

  (
    n1488_o2_n,
    n1488_o2
  );


  buf

  (
    n1602_o2_p,
    n1602_o2
  );


  not

  (
    n1602_o2_n,
    n1602_o2
  );


  buf

  (
    n517_o2_p,
    n517_o2
  );


  not

  (
    n517_o2_n,
    n517_o2
  );


  buf

  (
    n1603_o2_p,
    n1603_o2
  );


  not

  (
    n1603_o2_n,
    n1603_o2
  );


  buf

  (
    n509_o2_p,
    n509_o2
  );


  not

  (
    n509_o2_n,
    n509_o2
  );


  buf

  (
    n510_o2_p,
    n510_o2
  );


  not

  (
    n510_o2_n,
    n510_o2
  );


  buf

  (
    n579_o2_p,
    n579_o2
  );


  not

  (
    n579_o2_n,
    n579_o2
  );


  buf

  (
    n625_o2_p,
    n625_o2
  );


  not

  (
    n625_o2_n,
    n625_o2
  );


  buf

  (
    n679_o2_p,
    n679_o2
  );


  not

  (
    n679_o2_n,
    n679_o2
  );


  buf

  (
    n741_o2_p,
    n741_o2
  );


  not

  (
    n741_o2_n,
    n741_o2
  );


  buf

  (
    n811_o2_p,
    n811_o2
  );


  not

  (
    n811_o2_n,
    n811_o2
  );


  buf

  (
    n889_o2_p,
    n889_o2
  );


  not

  (
    n889_o2_n,
    n889_o2
  );


  buf

  (
    n975_o2_p,
    n975_o2
  );


  not

  (
    n975_o2_n,
    n975_o2
  );


  buf

  (
    n1069_o2_p,
    n1069_o2
  );


  not

  (
    n1069_o2_n,
    n1069_o2
  );


  buf

  (
    n1171_o2_p,
    n1171_o2
  );


  not

  (
    n1171_o2_n,
    n1171_o2
  );


  buf

  (
    n1281_o2_p,
    n1281_o2
  );


  not

  (
    n1281_o2_n,
    n1281_o2
  );


  buf

  (
    n1392_o2_p,
    n1392_o2
  );


  not

  (
    n1392_o2_n,
    n1392_o2
  );


  buf

  (
    n1501_o2_p,
    n1501_o2
  );


  not

  (
    n1501_o2_n,
    n1501_o2
  );


  buf

  (
    n541_o2_p,
    n541_o2
  );


  not

  (
    n541_o2_n,
    n541_o2
  );


  and

  (
    g389_p,
    n2491_lo_p,
    n2683_lo_p
  );


  or

  (
    g390_n,
    n3737_o2_p,
    n3736_o2_p
  );


  and

  (
    g391_p,
    n3801_o2_n,
    g390_n
  );


  and

  (
    g392_p,
    n3836_o2_p,
    n3885_o2_n
  );


  or

  (
    g393_n,
    n3902_o2_p,
    g392_p
  );


  and

  (
    g394_p,
    n4002_o2_p,
    n4052_o2_n
  );


  or

  (
    g395_n,
    n4067_o2_p,
    g394_p
  );


  and

  (
    g396_p,
    n4162_o2_p,
    n4212_o2_n
  );


  or

  (
    g397_n,
    n4227_o2_p,
    g396_p
  );


  and

  (
    g398_p,
    n4321_o2_p,
    n4367_o2_n
  );


  or

  (
    g399_n,
    n4383_o2_p,
    g398_p
  );


  and

  (
    g400_p,
    n4475_o2_p,
    n4523_o2_n
  );


  or

  (
    g401_n,
    n4537_o2_p,
    g400_p
  );


  and

  (
    g402_p,
    n4628_o2_p,
    n4674_o2_n
  );


  or

  (
    g403_n,
    n4688_o2_p,
    g402_p
  );


  and

  (
    g404_p,
    n4791_o2_p,
    n4835_o2_n
  );


  or

  (
    g405_n,
    n4868_o2_p,
    g404_p
  );


  and

  (
    g406_p,
    n5086_o2_p,
    n5130_o2_n
  );


  or

  (
    g407_n,
    n5188_o2_p,
    g406_p
  );


  and

  (
    g408_p,
    n5402_o2_p,
    n5445_o2_n
  );


  or

  (
    g409_n,
    n5500_o2_p,
    g408_p
  );


  and

  (
    g410_p,
    n5707_o2_p,
    n5745_o2_n
  );


  or

  (
    g411_n,
    n5801_o2_p,
    g410_p
  );


  and

  (
    g412_p,
    n6081_o2_p,
    n6120_o2_n
  );


  or

  (
    g413_n,
    n6203_o2_p,
    g412_p
  );


  and

  (
    g414_p,
    n6594_o2_p,
    n6631_o2_n
  );


  or

  (
    g415_n,
    n6725_o2_p,
    g414_p
  );


  and

  (
    g416_p,
    n1127_o2_p,
    n1231_o2_n
  );


  or

  (
    g417_n,
    n1232_o2_p,
    g416_p
  );


  and

  (
    g418_p,
    n1235_o2_p,
    n1347_o2_n
  );


  or

  (
    g419_n,
    n1348_o2_p,
    g418_p
  );


  or

  (
    g420_n,
    n1351_o2_p,
    n1461_o2_p
  );


  and

  (
    g421_p,
    n1463_o2_n,
    g420_n
  );


  and

  (
    g422_p,
    n1463_o2_p,
    n1573_o2_n
  );


  or

  (
    g423_n,
    n1574_o2_p,
    g422_p
  );


  and

  (
    g424_p,
    n1577_o2_p,
    n1678_o2_n
  );


  or

  (
    g425_n,
    n1679_o2_p,
    g424_p
  );


  and

  (
    g426_p,
    n1682_o2_p,
    n1775_o2_n
  );


  or

  (
    g427_n,
    n1776_o2_p,
    g426_p
  );


  and

  (
    g428_p,
    n1779_o2_p,
    n1864_o2_n
  );


  or

  (
    g429_n,
    n1865_o2_p,
    g428_p
  );


  and

  (
    g430_p,
    n1868_o2_p,
    n1945_o2_n
  );


  or

  (
    g431_n,
    n1946_o2_p_spl_,
    g430_p
  );


  and

  (
    g432_p,
    n1943_o2_p,
    n1946_o2_n
  );


  or

  (
    g432_n,
    n1943_o2_n,
    n1946_o2_p_spl_
  );


  and

  (
    g433_p,
    n2016_o2_p_spl_,
    n2017_o2_n
  );


  or

  (
    g433_n,
    n2016_o2_n_spl_,
    n2017_o2_p
  );


  and

  (
    g434_p,
    g432_n,
    g433_p
  );


  or

  (
    g434_n,
    g432_p_spl_,
    g433_n_spl_
  );


  and

  (
    g435_p,
    g432_p_spl_,
    g433_n_spl_
  );


  or

  (
    g436_n,
    g434_p_spl_,
    g435_p
  );


  and

  (
    g437_p,
    n2016_o2_p_spl_,
    g434_n
  );


  or

  (
    g437_n,
    n2016_o2_n_spl_,
    g434_p_spl_
  );


  and

  (
    g438_p,
    n2010_o2_p,
    n2013_o2_n
  );


  or

  (
    g438_n,
    n2010_o2_n,
    n2013_o2_p
  );


  and

  (
    g439_p,
    n2078_o2_n_spl_,
    n2079_o2_n
  );


  or

  (
    g439_n,
    n2078_o2_p_spl_,
    n2079_o2_p
  );


  and

  (
    g440_p,
    g438_n_spl_,
    g439_p_spl_
  );


  or

  (
    g440_n,
    g438_p_spl_,
    g439_n_spl_
  );


  and

  (
    g441_p,
    g438_p_spl_,
    g439_n_spl_
  );


  or

  (
    g441_n,
    g438_n_spl_,
    g439_p_spl_
  );


  and

  (
    g442_p,
    g440_n_spl_,
    g441_n
  );


  or

  (
    g442_n,
    g440_p_spl_,
    g441_p
  );


  and

  (
    g443_p,
    g437_n,
    g442_p
  );


  or

  (
    g443_n,
    g437_p_spl_,
    g442_n_spl_
  );


  and

  (
    g444_p,
    g437_p_spl_,
    g442_n_spl_
  );


  or

  (
    g445_n,
    g443_p_spl_,
    g444_p
  );


  and

  (
    g446_p,
    g440_n_spl_,
    g443_n
  );


  or

  (
    g446_n,
    g440_p_spl_,
    g443_p_spl_
  );


  and

  (
    g447_p,
    n2075_o2_p,
    n2078_o2_n_spl_
  );


  or

  (
    g447_n,
    n2075_o2_n,
    n2078_o2_p_spl_
  );


  and

  (
    g448_p,
    n2599_lo_p,
    n2863_lo_p_spl_00
  );


  or

  (
    g448_n,
    n2599_lo_n,
    n2863_lo_n_spl_00
  );


  and

  (
    g449_p,
    n2132_o2_p_spl_,
    n2133_o2_n
  );


  or

  (
    g449_n,
    n2132_o2_n_spl_,
    n2133_o2_p
  );


  and

  (
    g450_p,
    g448_n_spl_,
    g449_p_spl_
  );


  or

  (
    g450_n,
    g448_p_spl_,
    g449_n_spl_
  );


  and

  (
    g451_p,
    g448_p_spl_,
    g449_n_spl_
  );


  or

  (
    g451_n,
    g448_n_spl_,
    g449_p_spl_
  );


  and

  (
    g452_p,
    g450_n_spl_,
    g451_n
  );


  or

  (
    g452_n,
    g450_p_spl_,
    g451_p
  );


  and

  (
    g453_p,
    g447_n_spl_,
    g452_p_spl_
  );


  or

  (
    g453_n,
    g447_p_spl_,
    g452_n_spl_
  );


  and

  (
    g454_p,
    g447_p_spl_,
    g452_n_spl_
  );


  or

  (
    g454_n,
    g447_n_spl_,
    g452_p_spl_
  );


  and

  (
    g455_p,
    g453_n_spl_,
    g454_n
  );


  or

  (
    g455_n,
    g453_p_spl_,
    g454_p
  );


  and

  (
    g456_p,
    g446_n,
    g455_p
  );


  or

  (
    g456_n,
    g446_p_spl_,
    g455_n_spl_
  );


  and

  (
    g457_p,
    g446_p_spl_,
    g455_n_spl_
  );


  or

  (
    g458_n,
    g456_p_spl_,
    g457_p
  );


  and

  (
    g459_p,
    g453_n_spl_,
    g456_n
  );


  or

  (
    g459_n,
    g453_p_spl_,
    g456_p_spl_
  );


  and

  (
    g460_p,
    n2132_o2_p_spl_,
    g450_n_spl_
  );


  or

  (
    g460_n,
    n2132_o2_n_spl_,
    g450_p_spl_
  );


  and

  (
    g461_p,
    n2611_lo_p,
    n2863_lo_p_spl_00
  );


  or

  (
    g461_n,
    n2611_lo_n,
    n2863_lo_n_spl_00
  );


  and

  (
    g462_p,
    n2126_o2_p,
    n2129_o2_n
  );


  or

  (
    g462_n,
    n2126_o2_n,
    n2129_o2_p
  );


  and

  (
    g463_p,
    n2178_o2_n_spl_,
    n2179_o2_n
  );


  or

  (
    g463_n,
    n2178_o2_p_spl_,
    n2179_o2_p
  );


  and

  (
    g464_p,
    g462_n_spl_,
    g463_p_spl_
  );


  or

  (
    g464_n,
    g462_p_spl_,
    g463_n_spl_
  );


  and

  (
    g465_p,
    g462_p_spl_,
    g463_n_spl_
  );


  or

  (
    g465_n,
    g462_n_spl_,
    g463_p_spl_
  );


  and

  (
    g466_p,
    g464_n_spl_,
    g465_n
  );


  or

  (
    g466_n,
    g464_p_spl_,
    g465_p
  );


  and

  (
    g467_p,
    g461_n_spl_,
    g466_p_spl_
  );


  or

  (
    g467_n,
    g461_p_spl_,
    g466_n_spl_
  );


  and

  (
    g468_p,
    g461_p_spl_,
    g466_n_spl_
  );


  or

  (
    g468_n,
    g461_n_spl_,
    g466_p_spl_
  );


  and

  (
    g469_p,
    g467_n_spl_,
    g468_n
  );


  or

  (
    g469_n,
    g467_p_spl_,
    g468_p
  );


  and

  (
    g470_p,
    g460_n_spl_,
    g469_p_spl_
  );


  or

  (
    g470_n,
    g460_p_spl_,
    g469_n_spl_
  );


  and

  (
    g471_p,
    g460_p_spl_,
    g469_n_spl_
  );


  or

  (
    g471_n,
    g460_n_spl_,
    g469_p_spl_
  );


  and

  (
    g472_p,
    g470_n_spl_,
    g471_n
  );


  or

  (
    g472_n,
    g470_p_spl_,
    g471_p
  );


  and

  (
    g473_p,
    g459_n,
    g472_p
  );


  or

  (
    g473_n,
    g459_p_spl_,
    g472_n_spl_
  );


  and

  (
    g474_p,
    g459_p_spl_,
    g472_n_spl_
  );


  or

  (
    g475_n,
    g473_p_spl_,
    g474_p
  );


  and

  (
    g476_p,
    g470_n_spl_,
    g473_n
  );


  or

  (
    g476_n,
    g470_p_spl_,
    g473_p_spl_
  );


  and

  (
    g477_p,
    g464_n_spl_,
    g467_n_spl_
  );


  or

  (
    g477_n,
    g464_p_spl_,
    g467_p_spl_
  );


  and

  (
    g478_p,
    n2623_lo_p,
    n2863_lo_p_spl_01
  );


  or

  (
    g478_n,
    n2623_lo_n,
    n2863_lo_n_spl_01
  );


  and

  (
    g479_p,
    n2175_o2_p,
    n2178_o2_n_spl_
  );


  or

  (
    g479_n,
    n2175_o2_n,
    n2178_o2_p_spl_
  );


  and

  (
    g480_p,
    n2635_lo_p_spl_,
    n2851_lo_p_spl_0
  );


  or

  (
    g480_n,
    n2635_lo_n_spl_,
    n2851_lo_n_spl_0
  );


  and

  (
    g481_p,
    n2216_o2_p_spl_,
    n2217_o2_n
  );


  or

  (
    g481_n,
    n2216_o2_n_spl_,
    n2217_o2_p
  );


  and

  (
    g482_p,
    g480_n_spl_,
    g481_p_spl_
  );


  or

  (
    g482_n,
    g480_p_spl_,
    g481_n_spl_
  );


  and

  (
    g483_p,
    g480_p_spl_,
    g481_n_spl_
  );


  or

  (
    g483_n,
    g480_n_spl_,
    g481_p_spl_
  );


  and

  (
    g484_p,
    g482_n_spl_,
    g483_n
  );


  or

  (
    g484_n,
    g482_p_spl_,
    g483_p
  );


  and

  (
    g485_p,
    g479_n_spl_,
    g484_p_spl_
  );


  or

  (
    g485_n,
    g479_p_spl_,
    g484_n_spl_
  );


  and

  (
    g486_p,
    g479_p_spl_,
    g484_n_spl_
  );


  or

  (
    g486_n,
    g479_n_spl_,
    g484_p_spl_
  );


  and

  (
    g487_p,
    g485_n_spl_,
    g486_n
  );


  or

  (
    g487_n,
    g485_p_spl_,
    g486_p
  );


  and

  (
    g488_p,
    g478_n_spl_,
    g487_p_spl_
  );


  or

  (
    g488_n,
    g478_p_spl_,
    g487_n_spl_
  );


  and

  (
    g489_p,
    g478_p_spl_,
    g487_n_spl_
  );


  or

  (
    g489_n,
    g478_n_spl_,
    g487_p_spl_
  );


  and

  (
    g490_p,
    g488_n_spl_,
    g489_n
  );


  or

  (
    g490_n,
    g488_p_spl_,
    g489_p
  );


  and

  (
    g491_p,
    g477_n_spl_,
    g490_p_spl_
  );


  or

  (
    g491_n,
    g477_p_spl_,
    g490_n_spl_
  );


  and

  (
    g492_p,
    g477_p_spl_,
    g490_n_spl_
  );


  or

  (
    g492_n,
    g477_n_spl_,
    g490_p_spl_
  );


  and

  (
    g493_p,
    g491_n_spl_,
    g492_n
  );


  or

  (
    g493_n,
    g491_p_spl_,
    g492_p
  );


  and

  (
    g494_p,
    g476_n,
    g493_p
  );


  or

  (
    g494_n,
    g476_p_spl_,
    g493_n_spl_
  );


  and

  (
    g495_p,
    g476_p_spl_,
    g493_n_spl_
  );


  or

  (
    g496_n,
    g494_p_spl_,
    g495_p
  );


  and

  (
    g497_p,
    g491_n_spl_,
    g494_n
  );


  or

  (
    g497_n,
    g491_p_spl_,
    g494_p_spl_
  );


  and

  (
    g498_p,
    g485_n_spl_,
    g488_n_spl_
  );


  or

  (
    g498_n,
    g485_p_spl_,
    g488_p_spl_
  );


  and

  (
    g499_p,
    n2635_lo_p_spl_,
    n2863_lo_p_spl_01
  );


  or

  (
    g499_n,
    n2635_lo_n_spl_,
    n2863_lo_n_spl_01
  );


  and

  (
    g500_p,
    n2216_o2_p_spl_,
    g482_n_spl_
  );


  or

  (
    g500_n,
    n2216_o2_n_spl_,
    g482_p_spl_
  );


  and

  (
    g501_p,
    n2647_lo_p_spl_,
    n2851_lo_p_spl_0
  );


  or

  (
    g501_n,
    n2647_lo_n_spl_,
    n2851_lo_n_spl_0
  );


  and

  (
    g502_p,
    n2210_o2_p,
    n2213_o2_n
  );


  or

  (
    g502_n,
    n2210_o2_n,
    n2213_o2_p
  );


  and

  (
    g503_p,
    n2246_o2_n_spl_,
    n2247_o2_n
  );


  or

  (
    g503_n,
    n2246_o2_p_spl_,
    n2247_o2_p
  );


  and

  (
    g504_p,
    g502_n_spl_,
    g503_p_spl_
  );


  or

  (
    g504_n,
    g502_p_spl_,
    g503_n_spl_
  );


  and

  (
    g505_p,
    g502_p_spl_,
    g503_n_spl_
  );


  or

  (
    g505_n,
    g502_n_spl_,
    g503_p_spl_
  );


  and

  (
    g506_p,
    g504_n_spl_,
    g505_n
  );


  or

  (
    g506_n,
    g504_p_spl_,
    g505_p
  );


  and

  (
    g507_p,
    g501_n_spl_,
    g506_p_spl_
  );


  or

  (
    g507_n,
    g501_p_spl_,
    g506_n_spl_
  );


  and

  (
    g508_p,
    g501_p_spl_,
    g506_n_spl_
  );


  or

  (
    g508_n,
    g501_n_spl_,
    g506_p_spl_
  );


  and

  (
    g509_p,
    g507_n_spl_,
    g508_n
  );


  or

  (
    g509_n,
    g507_p_spl_,
    g508_p
  );


  and

  (
    g510_p,
    g500_n_spl_,
    g509_p_spl_
  );


  or

  (
    g510_n,
    g500_p_spl_,
    g509_n_spl_
  );


  and

  (
    g511_p,
    g500_p_spl_,
    g509_n_spl_
  );


  or

  (
    g511_n,
    g500_n_spl_,
    g509_p_spl_
  );


  and

  (
    g512_p,
    g510_n_spl_,
    g511_n
  );


  or

  (
    g512_n,
    g510_p_spl_,
    g511_p
  );


  and

  (
    g513_p,
    g499_n_spl_,
    g512_p_spl_
  );


  or

  (
    g513_n,
    g499_p_spl_,
    g512_n_spl_
  );


  and

  (
    g514_p,
    g499_p_spl_,
    g512_n_spl_
  );


  or

  (
    g514_n,
    g499_n_spl_,
    g512_p_spl_
  );


  and

  (
    g515_p,
    g513_n_spl_,
    g514_n
  );


  or

  (
    g515_n,
    g513_p_spl_,
    g514_p
  );


  and

  (
    g516_p,
    g498_n_spl_,
    g515_p_spl_
  );


  or

  (
    g516_n,
    g498_p_spl_,
    g515_n_spl_
  );


  and

  (
    g517_p,
    g498_p_spl_,
    g515_n_spl_
  );


  or

  (
    g517_n,
    g498_n_spl_,
    g515_p_spl_
  );


  and

  (
    g518_p,
    g516_n_spl_,
    g517_n
  );


  or

  (
    g518_n,
    g516_p_spl_,
    g517_p
  );


  and

  (
    g519_p,
    g497_n,
    g518_p
  );


  or

  (
    g519_n,
    g497_p_spl_,
    g518_n_spl_
  );


  and

  (
    g520_p,
    g497_p_spl_,
    g518_n_spl_
  );


  or

  (
    g521_n,
    g519_p_spl_,
    g520_p
  );


  and

  (
    g522_p,
    g516_n_spl_,
    g519_n
  );


  or

  (
    g522_n,
    g516_p_spl_,
    g519_p_spl_
  );


  and

  (
    g523_p,
    g510_n_spl_,
    g513_n_spl_
  );


  or

  (
    g523_n,
    g510_p_spl_,
    g513_p_spl_
  );


  and

  (
    g524_p,
    n2647_lo_p_spl_,
    n2863_lo_p_spl_10
  );


  or

  (
    g524_n,
    n2647_lo_n_spl_,
    n2863_lo_n_spl_10
  );


  and

  (
    g525_p,
    g504_n_spl_,
    g507_n_spl_
  );


  or

  (
    g525_n,
    g504_p_spl_,
    g507_p_spl_
  );


  and

  (
    g526_p,
    n2659_lo_p_spl_,
    n2851_lo_p_spl_1
  );


  or

  (
    g526_n,
    n2659_lo_n_spl_,
    n2851_lo_n_spl_1
  );


  and

  (
    g527_p,
    n2671_lo_p_spl_0,
    n2839_lo_p
  );


  or

  (
    g527_n,
    n2671_lo_n_spl_0,
    n2839_lo_n
  );


  and

  (
    g528_p,
    n2243_o2_p,
    n2246_o2_n_spl_
  );


  or

  (
    g528_n,
    n2243_o2_n,
    n2246_o2_p_spl_
  );


  and

  (
    g529_p,
    g527_n_spl_,
    g528_n_spl_
  );


  or

  (
    g529_n,
    g527_p_spl_,
    g528_p_spl_
  );


  and

  (
    g530_p,
    g527_p_spl_,
    g528_p_spl_
  );


  or

  (
    g530_n,
    g527_n_spl_,
    g528_n_spl_
  );


  and

  (
    g531_p,
    g529_n_spl_,
    g530_n
  );


  or

  (
    g531_n,
    g529_p_spl_,
    g530_p
  );


  and

  (
    g532_p,
    g526_n_spl_,
    g531_p_spl_
  );


  or

  (
    g532_n,
    g526_p_spl_,
    g531_n_spl_
  );


  and

  (
    g533_p,
    g526_p_spl_,
    g531_n_spl_
  );


  or

  (
    g533_n,
    g526_n_spl_,
    g531_p_spl_
  );


  and

  (
    g534_p,
    g532_n_spl_,
    g533_n
  );


  or

  (
    g534_n,
    g532_p_spl_,
    g533_p
  );


  and

  (
    g535_p,
    g525_n_spl_,
    g534_p_spl_
  );


  or

  (
    g535_n,
    g525_p_spl_,
    g534_n_spl_
  );


  and

  (
    g536_p,
    g525_p_spl_,
    g534_n_spl_
  );


  or

  (
    g536_n,
    g525_n_spl_,
    g534_p_spl_
  );


  and

  (
    g537_p,
    g535_n_spl_,
    g536_n
  );


  or

  (
    g537_n,
    g535_p_spl_,
    g536_p
  );


  and

  (
    g538_p,
    g524_n_spl_,
    g537_p_spl_
  );


  or

  (
    g538_n,
    g524_p_spl_,
    g537_n_spl_
  );


  and

  (
    g539_p,
    g524_p_spl_,
    g537_n_spl_
  );


  or

  (
    g539_n,
    g524_n_spl_,
    g537_p_spl_
  );


  and

  (
    g540_p,
    g538_n_spl_,
    g539_n
  );


  or

  (
    g540_n,
    g538_p_spl_,
    g539_p
  );


  and

  (
    g541_p,
    g523_n_spl_,
    g540_p_spl_
  );


  or

  (
    g541_n,
    g523_p_spl_,
    g540_n_spl_
  );


  and

  (
    g542_p,
    g523_p_spl_,
    g540_n_spl_
  );


  or

  (
    g542_n,
    g523_n_spl_,
    g540_p_spl_
  );


  and

  (
    g543_p,
    g541_n_spl_,
    g542_n
  );


  or

  (
    g543_n,
    g541_p_spl_,
    g542_p
  );


  and

  (
    g544_p,
    g522_n,
    g543_p
  );


  or

  (
    g544_n,
    g522_p_spl_,
    g543_n_spl_
  );


  and

  (
    g545_p,
    g522_p_spl_,
    g543_n_spl_
  );


  or

  (
    g546_n,
    g544_p_spl_,
    g545_p
  );


  and

  (
    g547_p,
    g541_n_spl_,
    g544_n
  );


  or

  (
    g547_n,
    g541_p_spl_,
    g544_p_spl_
  );


  and

  (
    g548_p,
    g535_n_spl_,
    g538_n_spl_
  );


  or

  (
    g548_n,
    g535_p_spl_,
    g538_p_spl_
  );


  and

  (
    g549_p,
    n2659_lo_p_spl_,
    n2863_lo_p_spl_10
  );


  or

  (
    g549_n,
    n2659_lo_n_spl_,
    n2863_lo_n_spl_10
  );


  and

  (
    g550_p,
    n2671_lo_p_spl_0,
    n2851_lo_p_spl_1
  );


  or

  (
    g550_n,
    n2671_lo_n_spl_0,
    n2851_lo_n_spl_1
  );


  and

  (
    g551_p,
    g529_n_spl_,
    g532_n_spl_
  );


  or

  (
    g551_n,
    g529_p_spl_,
    g532_p_spl_
  );


  and

  (
    g552_p,
    g550_n_spl_,
    g551_n_spl_
  );


  or

  (
    g552_n,
    g550_p_spl_,
    g551_p_spl_
  );


  and

  (
    g553_p,
    g550_p_spl_,
    g551_p_spl_
  );


  or

  (
    g553_n,
    g550_n_spl_,
    g551_n_spl_
  );


  and

  (
    g554_p,
    g552_n_spl_,
    g553_n
  );


  or

  (
    g554_n,
    g552_p_spl_,
    g553_p
  );


  and

  (
    g555_p,
    g549_n_spl_,
    g554_p_spl_
  );


  or

  (
    g555_n,
    g549_p_spl_,
    g554_n_spl_
  );


  and

  (
    g556_p,
    g549_p_spl_,
    g554_n_spl_
  );


  or

  (
    g556_n,
    g549_n_spl_,
    g554_p_spl_
  );


  and

  (
    g557_p,
    g555_n_spl_,
    g556_n
  );


  or

  (
    g557_n,
    g555_p_spl_,
    g556_p
  );


  and

  (
    g558_p,
    g548_n_spl_,
    g557_p_spl_
  );


  or

  (
    g558_n,
    g548_p_spl_,
    g557_n_spl_
  );


  and

  (
    g559_p,
    g548_p_spl_,
    g557_n_spl_
  );


  or

  (
    g559_n,
    g548_n_spl_,
    g557_p_spl_
  );


  and

  (
    g560_p,
    g558_n_spl_,
    g559_n
  );


  or

  (
    g560_n,
    g558_p_spl_,
    g559_p
  );


  and

  (
    g561_p,
    g547_n,
    g560_p
  );


  or

  (
    g561_n,
    g547_p_spl_,
    g560_n_spl_
  );


  and

  (
    g562_p,
    g547_p_spl_,
    g560_n_spl_
  );


  or

  (
    g563_n,
    g561_p_spl_,
    g562_p
  );


  and

  (
    g564_p,
    n2671_lo_p_spl_,
    n2863_lo_p_spl_1
  );


  or

  (
    g564_n,
    n2671_lo_n_spl_,
    n2863_lo_n_spl_1
  );


  and

  (
    g565_p,
    g552_n_spl_,
    g555_n_spl_
  );


  or

  (
    g565_n,
    g552_p_spl_,
    g555_p_spl_
  );


  and

  (
    g566_p,
    g564_n_spl_,
    g565_n_spl_
  );


  or

  (
    g566_n,
    g564_p_spl_,
    g565_p_spl_
  );


  and

  (
    g567_p,
    g558_n_spl_,
    g561_n
  );


  or

  (
    g567_n,
    g558_p_spl_,
    g561_p_spl_
  );


  and

  (
    g568_p,
    g564_p_spl_,
    g565_p_spl_
  );


  or

  (
    g568_n,
    g564_n_spl_,
    g565_n_spl_
  );


  and

  (
    g569_p,
    g566_n_spl_,
    g568_n
  );


  or

  (
    g569_n,
    g566_p,
    g568_p
  );


  or

  (
    g570_n,
    g567_p,
    g569_n
  );


  and

  (
    g571_p,
    g566_n_spl_,
    g570_n_spl_
  );


  or

  (
    g572_n,
    g567_n,
    g569_p
  );


  and

  (
    g573_p,
    g570_n_spl_,
    g572_n
  );


  and

  (
    g574_p,
    n2848_lo_p_spl_000,
    n4908_o2_p_spl_
  );


  or

  (
    g574_n,
    n2848_lo_n_spl_000,
    n4908_o2_n_spl_
  );


  and

  (
    g575_p,
    n1121_o2_p,
    n1124_o2_n
  );


  or

  (
    g575_n,
    n1121_o2_n,
    n1124_o2_p_spl_
  );


  and

  (
    g576_p,
    n1226_o2_n,
    n1227_o2_n
  );


  or

  (
    g576_n,
    n1226_o2_p,
    n1227_o2_p
  );


  and

  (
    g577_p,
    g575_n_spl_,
    g576_p_spl_
  );


  or

  (
    g577_n,
    g575_p_spl_,
    g576_n_spl_
  );


  and

  (
    g578_p,
    g575_p_spl_,
    g576_n_spl_
  );


  or

  (
    g578_n,
    g575_n_spl_,
    g576_p_spl_
  );


  and

  (
    g579_p,
    g577_n_spl_,
    g578_n
  );


  or

  (
    g579_n,
    g577_p_spl_,
    g578_p
  );


  and

  (
    g580_p,
    g574_n,
    g579_p_spl_
  );


  or

  (
    g580_n,
    g574_p_spl_,
    g579_n
  );


  or

  (
    g581_n,
    n2860_lo_n_spl_000,
    n4908_o2_n_spl_
  );


  and

  (
    g582_p,
    g577_n_spl_,
    g580_n
  );


  or

  (
    g582_n,
    g577_p_spl_,
    g580_p_spl_
  );


  and

  (
    g583_p,
    n2848_lo_p_spl_000,
    n4867_o2_p_spl_
  );


  or

  (
    g583_n,
    n2848_lo_n_spl_000,
    n4867_o2_n_spl_
  );


  and

  (
    g584_p,
    n1238_o2_n_spl_,
    n1338_o2_n_spl_
  );


  or

  (
    g584_n,
    n1238_o2_p_spl_,
    n1338_o2_p_spl_
  );


  and

  (
    g585_p,
    n1238_o2_p_spl_,
    n1338_o2_p_spl_
  );


  or

  (
    g585_n,
    n1238_o2_n_spl_,
    n1338_o2_n_spl_
  );


  and

  (
    g586_p,
    g584_n_spl_,
    g585_n
  );


  or

  (
    g586_n,
    g584_p_spl_,
    g585_p
  );


  and

  (
    g587_p,
    g583_n_spl_,
    g586_p_spl_
  );


  or

  (
    g587_n,
    g583_p_spl_,
    g586_n_spl_
  );


  and

  (
    g588_p,
    g583_p_spl_,
    g586_n_spl_
  );


  or

  (
    g588_n,
    g583_n_spl_,
    g586_p_spl_
  );


  and

  (
    g589_p,
    g587_n_spl_,
    g588_n
  );


  or

  (
    g589_n,
    g587_p_spl_,
    g588_p
  );


  and

  (
    g590_p,
    g582_n_spl_,
    g589_p_spl_
  );


  or

  (
    g590_n,
    g582_p,
    g589_n
  );


  or

  (
    g591_n,
    g582_n_spl_,
    g589_p_spl_
  );


  and

  (
    g592_p,
    g590_n,
    g591_n
  );


  and

  (
    g593_p,
    g581_n_spl_,
    g592_p_spl_
  );


  or

  (
    g594_n,
    g590_p,
    g593_p_spl_
  );


  and

  (
    g595_p,
    n2860_lo_p_spl_00,
    n4867_o2_p_spl_
  );


  or

  (
    g595_n,
    n2860_lo_n_spl_000,
    n4867_o2_n_spl_
  );


  and

  (
    g596_p,
    g584_n_spl_,
    g587_n_spl_
  );


  or

  (
    g596_n,
    g584_p_spl_,
    g587_p_spl_
  );


  and

  (
    g597_p,
    n2848_lo_p_spl_001,
    n4836_o2_p_spl_
  );


  or

  (
    g597_n,
    n2848_lo_n_spl_001,
    n4836_o2_n_spl_
  );


  and

  (
    g598_p,
    n1355_o2_n_spl_,
    n1449_o2_n_spl_
  );


  or

  (
    g598_n,
    n1355_o2_p_spl_,
    n1449_o2_p_spl_
  );


  and

  (
    g599_p,
    n1355_o2_p_spl_,
    n1449_o2_p_spl_
  );


  or

  (
    g599_n,
    n1355_o2_n_spl_,
    n1449_o2_n_spl_
  );


  and

  (
    g600_p,
    g598_n_spl_,
    g599_n
  );


  or

  (
    g600_n,
    g598_p_spl_,
    g599_p
  );


  and

  (
    g601_p,
    g597_n_spl_,
    g600_p_spl_
  );


  or

  (
    g601_n,
    g597_p_spl_,
    g600_n_spl_
  );


  and

  (
    g602_p,
    g597_p_spl_,
    g600_n_spl_
  );


  or

  (
    g602_n,
    g597_n_spl_,
    g600_p_spl_
  );


  and

  (
    g603_p,
    g601_n_spl_,
    g602_n
  );


  or

  (
    g603_n,
    g601_p_spl_,
    g602_p
  );


  and

  (
    g604_p,
    g596_n_spl_,
    g603_p_spl_
  );


  or

  (
    g604_n,
    g596_p_spl_,
    g603_n_spl_
  );


  and

  (
    g605_p,
    g596_p_spl_,
    g603_n_spl_
  );


  or

  (
    g605_n,
    g596_n_spl_,
    g603_p_spl_
  );


  and

  (
    g606_p,
    g604_n_spl_,
    g605_n
  );


  or

  (
    g606_n,
    g604_p_spl_,
    g605_p
  );


  and

  (
    g607_p,
    g595_n_spl_,
    g606_p_spl_
  );


  or

  (
    g607_n,
    g595_p,
    g606_n
  );


  or

  (
    g608_n,
    g595_n_spl_,
    g606_p_spl_
  );


  and

  (
    g609_p,
    g607_n_spl_,
    g608_n
  );


  or

  (
    g610_n,
    g594_n_spl_,
    g609_p_spl_
  );


  and

  (
    g611_p,
    g604_n_spl_,
    g607_n_spl_
  );


  or

  (
    g611_n,
    g604_p_spl_,
    g607_p
  );


  and

  (
    g612_p,
    n2860_lo_p_spl_00,
    n4836_o2_p_spl_
  );


  or

  (
    g612_n,
    n2860_lo_n_spl_00,
    n4836_o2_n_spl_
  );


  and

  (
    g613_p,
    g598_n_spl_,
    g601_n_spl_
  );


  or

  (
    g613_n,
    g598_p_spl_,
    g601_p_spl_
  );


  and

  (
    g614_p,
    n2848_lo_p_spl_001,
    n4837_o2_p_spl_
  );


  or

  (
    g614_n,
    n2848_lo_n_spl_001,
    n4837_o2_n_spl_
  );


  and

  (
    g615_p,
    n1469_o2_n_spl_,
    n1558_o2_n_spl_
  );


  or

  (
    g615_n,
    n1469_o2_p_spl_,
    n1558_o2_p_spl_
  );


  and

  (
    g616_p,
    n1469_o2_p_spl_,
    n1558_o2_p_spl_
  );


  or

  (
    g616_n,
    n1469_o2_n_spl_,
    n1558_o2_n_spl_
  );


  and

  (
    g617_p,
    g615_n_spl_,
    g616_n
  );


  or

  (
    g617_n,
    g615_p_spl_,
    g616_p
  );


  and

  (
    g618_p,
    g614_n_spl_,
    g617_p_spl_
  );


  or

  (
    g618_n,
    g614_p_spl_,
    g617_n_spl_
  );


  and

  (
    g619_p,
    g614_p_spl_,
    g617_n_spl_
  );


  or

  (
    g619_n,
    g614_n_spl_,
    g617_p_spl_
  );


  and

  (
    g620_p,
    g618_n_spl_,
    g619_n
  );


  or

  (
    g620_n,
    g618_p_spl_,
    g619_p
  );


  and

  (
    g621_p,
    g613_n_spl_,
    g620_p_spl_
  );


  or

  (
    g621_n,
    g613_p_spl_,
    g620_n_spl_
  );


  and

  (
    g622_p,
    g613_p_spl_,
    g620_n_spl_
  );


  or

  (
    g622_n,
    g613_n_spl_,
    g620_p_spl_
  );


  and

  (
    g623_p,
    g621_n_spl_,
    g622_n
  );


  or

  (
    g623_n,
    g621_p_spl_,
    g622_p
  );


  and

  (
    g624_p,
    g612_n_spl_,
    g623_p_spl_
  );


  or

  (
    g624_n,
    g612_p_spl_,
    g623_n_spl_
  );


  and

  (
    g625_p,
    g612_p_spl_,
    g623_n_spl_
  );


  or

  (
    g625_n,
    g612_n_spl_,
    g623_p_spl_
  );


  and

  (
    g626_p,
    g624_n_spl_,
    g625_n
  );


  or

  (
    g626_n,
    g624_p_spl_,
    g625_p
  );


  and

  (
    g627_p,
    g611_n_spl_,
    g626_p_spl_
  );


  or

  (
    g627_n,
    g611_p,
    g626_n
  );


  or

  (
    g628_n,
    g611_n_spl_,
    g626_p_spl_
  );


  and

  (
    g629_p,
    g627_n,
    g628_n
  );


  and

  (
    g630_p,
    n6148_o2_p_spl_00,
    lo102_buf_o2_p_spl_000
  );


  or

  (
    g630_n,
    n6148_o2_n_spl_00,
    lo102_buf_o2_n_spl_000
  );


  and

  (
    g631_p,
    g610_n_spl_,
    g629_p_spl_
  );


  and

  (
    g632_p,
    n708_o2_n_spl_,
    n768_o2_n_spl_
  );


  or

  (
    g632_n,
    n708_o2_p_spl_,
    n768_o2_p_spl_
  );


  and

  (
    g633_p,
    n708_o2_p_spl_,
    n768_o2_p_spl_
  );


  or

  (
    g633_n,
    n708_o2_n_spl_,
    n768_o2_n_spl_
  );


  and

  (
    g634_p,
    g632_n_spl_,
    g633_n
  );


  or

  (
    g634_n,
    g632_p_spl_,
    g633_p
  );


  and

  (
    g635_p,
    g630_n,
    g634_p_spl_
  );


  or

  (
    g635_n,
    g630_p_spl_,
    g634_n
  );


  or

  (
    g636_n,
    g627_p,
    g631_p_spl_
  );


  and

  (
    g637_p,
    g621_n_spl_,
    g624_n_spl_
  );


  or

  (
    g637_n,
    g621_p_spl_,
    g624_p_spl_
  );


  and

  (
    g638_p,
    n2860_lo_p_spl_01,
    n4837_o2_p_spl_
  );


  or

  (
    g638_n,
    n2860_lo_n_spl_01,
    n4837_o2_n_spl_
  );


  and

  (
    g639_p,
    g615_n_spl_,
    g618_n_spl_
  );


  or

  (
    g639_n,
    g615_p_spl_,
    g618_p_spl_
  );


  and

  (
    g640_p,
    n2848_lo_p_spl_010,
    n4838_o2_p_spl_
  );


  or

  (
    g640_n,
    n2848_lo_n_spl_010,
    n4838_o2_n_spl_
  );


  and

  (
    g641_p,
    n1553_o2_p,
    n1556_o2_n
  );


  or

  (
    g641_n,
    n1553_o2_n,
    n1556_o2_p
  );


  and

  (
    g642_p,
    n1583_o2_n_spl_,
    n1660_o2_p_spl_
  );


  or

  (
    g642_n,
    n1583_o2_p_spl_,
    n1660_o2_n_spl_
  );


  and

  (
    g643_p,
    n1583_o2_p_spl_,
    n1660_o2_n_spl_
  );


  or

  (
    g643_n,
    n1583_o2_n_spl_,
    n1660_o2_p_spl_
  );


  and

  (
    g644_p,
    g642_n_spl_,
    g643_n
  );


  or

  (
    g644_n,
    g642_p_spl_,
    g643_p
  );


  and

  (
    g645_p,
    g641_n_spl_,
    g644_p_spl_
  );


  or

  (
    g645_n,
    g641_p_spl_,
    g644_n_spl_
  );


  and

  (
    g646_p,
    g641_p_spl_,
    g644_n_spl_
  );


  or

  (
    g646_n,
    g641_n_spl_,
    g644_p_spl_
  );


  and

  (
    g647_p,
    g645_n_spl_,
    g646_n
  );


  or

  (
    g647_n,
    g645_p_spl_,
    g646_p
  );


  and

  (
    g648_p,
    g640_n_spl_,
    g647_p_spl_
  );


  or

  (
    g648_n,
    g640_p_spl_,
    g647_n_spl_
  );


  and

  (
    g649_p,
    g640_p_spl_,
    g647_n_spl_
  );


  or

  (
    g649_n,
    g640_n_spl_,
    g647_p_spl_
  );


  and

  (
    g650_p,
    g648_n_spl_,
    g649_n
  );


  or

  (
    g650_n,
    g648_p_spl_,
    g649_p
  );


  and

  (
    g651_p,
    g639_n_spl_,
    g650_p_spl_
  );


  or

  (
    g651_n,
    g639_p_spl_,
    g650_n_spl_
  );


  and

  (
    g652_p,
    g639_p_spl_,
    g650_n_spl_
  );


  or

  (
    g652_n,
    g639_n_spl_,
    g650_p_spl_
  );


  and

  (
    g653_p,
    g651_n_spl_,
    g652_n
  );


  or

  (
    g653_n,
    g651_p_spl_,
    g652_p
  );


  and

  (
    g654_p,
    g638_n_spl_,
    g653_p_spl_
  );


  or

  (
    g654_n,
    g638_p_spl_,
    g653_n_spl_
  );


  and

  (
    g655_p,
    g638_p_spl_,
    g653_n_spl_
  );


  or

  (
    g655_n,
    g638_n_spl_,
    g653_p_spl_
  );


  and

  (
    g656_p,
    g654_n_spl_,
    g655_n
  );


  or

  (
    g656_n,
    g654_p_spl_,
    g655_p
  );


  and

  (
    g657_p,
    g637_n_spl_,
    g656_p_spl_
  );


  or

  (
    g657_n,
    g637_p,
    g656_n
  );


  or

  (
    g658_n,
    g637_n_spl_,
    g656_p_spl_
  );


  and

  (
    g659_p,
    g657_n,
    g658_n
  );


  and

  (
    g660_p,
    n2797_lo_p_spl_000,
    n6148_o2_p_spl_00
  );


  or

  (
    g660_n,
    n2797_lo_n_spl_000,
    n6148_o2_n_spl_00
  );


  and

  (
    g661_p,
    g636_n_spl_,
    g659_p_spl_
  );


  and

  (
    g662_p,
    g632_n_spl_,
    g635_n
  );


  or

  (
    g662_n,
    g632_p_spl_,
    g635_p_spl_
  );


  and

  (
    g663_p,
    n6053_o2_p_spl_00,
    lo102_buf_o2_p_spl_000
  );


  or

  (
    g663_n,
    n6053_o2_n_spl_00,
    lo102_buf_o2_n_spl_000
  );


  and

  (
    g664_p,
    n839_o2_p_spl_,
    n840_o2_n
  );


  or

  (
    g664_n,
    n839_o2_n_spl_,
    n840_o2_p
  );


  and

  (
    g665_p,
    g663_n_spl_,
    g664_p_spl_
  );


  or

  (
    g665_n,
    g663_p_spl_,
    g664_n_spl_
  );


  and

  (
    g666_p,
    g663_p_spl_,
    g664_n_spl_
  );


  or

  (
    g666_n,
    g663_n_spl_,
    g664_p_spl_
  );


  and

  (
    g667_p,
    g665_n_spl_,
    g666_n
  );


  or

  (
    g667_n,
    g665_p_spl_,
    g666_p
  );


  and

  (
    g668_p,
    g662_n_spl_,
    g667_p_spl_
  );


  or

  (
    g668_n,
    g662_p_spl_,
    g667_n_spl_
  );


  and

  (
    g669_p,
    g662_p_spl_,
    g667_n_spl_
  );


  or

  (
    g669_n,
    g662_n_spl_,
    g667_p_spl_
  );


  and

  (
    g670_p,
    g668_n_spl_,
    g669_n
  );


  or

  (
    g670_n,
    g668_p_spl_,
    g669_p
  );


  and

  (
    g671_p,
    g660_n,
    g670_p_spl_
  );


  or

  (
    g671_n,
    g660_p_spl_,
    g670_n
  );


  and

  (
    g672_p,
    lo002_buf_o2_p_spl_00,
    lo082_buf_o2_p_spl_0
  );


  or

  (
    g672_n,
    lo002_buf_o2_n_spl_00,
    lo082_buf_o2_n_spl_0
  );


  and

  (
    g673_p,
    n509_o2_p_spl_,
    n510_o2_n
  );


  or

  (
    g673_n,
    n509_o2_n_spl_,
    n510_o2_p
  );


  or

  (
    g674_n,
    g657_p,
    g661_p_spl_
  );


  and

  (
    g675_p,
    g651_n_spl_,
    g654_n_spl_
  );


  or

  (
    g675_n,
    g651_p_spl_,
    g654_p_spl_
  );


  and

  (
    g676_p,
    n2860_lo_p_spl_01,
    n4838_o2_p_spl_
  );


  or

  (
    g676_n,
    n2860_lo_n_spl_01,
    n4838_o2_n_spl_
  );


  and

  (
    g677_p,
    g645_n_spl_,
    g648_n_spl_
  );


  or

  (
    g677_n,
    g645_p_spl_,
    g648_p_spl_
  );


  and

  (
    g678_p,
    n2848_lo_p_spl_010,
    n4839_o2_p_spl_
  );


  or

  (
    g678_n,
    n2848_lo_n_spl_010,
    n4839_o2_n_spl_
  );


  and

  (
    g679_p,
    n1658_o2_p,
    g642_n_spl_
  );


  or

  (
    g679_n,
    n1658_o2_n,
    g642_p_spl_
  );


  and

  (
    g680_p,
    n4840_o2_p_spl_0,
    lo118_buf_o2_p_spl_000
  );


  or

  (
    g680_n,
    n4840_o2_n_spl_0,
    lo118_buf_o2_n_spl_000
  );


  and

  (
    g681_p,
    n1689_o2_n_spl_,
    n1754_o2_n_spl_
  );


  or

  (
    g681_n,
    n1689_o2_p_spl_,
    n1754_o2_p_spl_
  );


  and

  (
    g682_p,
    n1689_o2_p_spl_,
    n1754_o2_p_spl_
  );


  or

  (
    g682_n,
    n1689_o2_n_spl_,
    n1754_o2_n_spl_
  );


  and

  (
    g683_p,
    g681_n_spl_,
    g682_n
  );


  or

  (
    g683_n,
    g681_p_spl_,
    g682_p
  );


  and

  (
    g684_p,
    g680_n_spl_,
    g683_p_spl_
  );


  or

  (
    g684_n,
    g680_p_spl_,
    g683_n_spl_
  );


  and

  (
    g685_p,
    g680_p_spl_,
    g683_n_spl_
  );


  or

  (
    g685_n,
    g680_n_spl_,
    g683_p_spl_
  );


  and

  (
    g686_p,
    g684_n_spl_,
    g685_n
  );


  or

  (
    g686_n,
    g684_p_spl_,
    g685_p
  );


  and

  (
    g687_p,
    g679_n_spl_,
    g686_p_spl_
  );


  or

  (
    g687_n,
    g679_p_spl_,
    g686_n_spl_
  );


  and

  (
    g688_p,
    g679_p_spl_,
    g686_n_spl_
  );


  or

  (
    g688_n,
    g679_n_spl_,
    g686_p_spl_
  );


  and

  (
    g689_p,
    g687_n_spl_,
    g688_n
  );


  or

  (
    g689_n,
    g687_p_spl_,
    g688_p
  );


  and

  (
    g690_p,
    g678_n_spl_,
    g689_p_spl_
  );


  or

  (
    g690_n,
    g678_p_spl_,
    g689_n_spl_
  );


  and

  (
    g691_p,
    g678_p_spl_,
    g689_n_spl_
  );


  or

  (
    g691_n,
    g678_n_spl_,
    g689_p_spl_
  );


  and

  (
    g692_p,
    g690_n_spl_,
    g691_n
  );


  or

  (
    g692_n,
    g690_p_spl_,
    g691_p
  );


  and

  (
    g693_p,
    g677_n_spl_,
    g692_p_spl_
  );


  or

  (
    g693_n,
    g677_p_spl_,
    g692_n_spl_
  );


  and

  (
    g694_p,
    g677_p_spl_,
    g692_n_spl_
  );


  or

  (
    g694_n,
    g677_n_spl_,
    g692_p_spl_
  );


  and

  (
    g695_p,
    g693_n_spl_,
    g694_n
  );


  or

  (
    g695_n,
    g693_p_spl_,
    g694_p
  );


  and

  (
    g696_p,
    g676_n_spl_,
    g695_p_spl_
  );


  or

  (
    g696_n,
    g676_p_spl_,
    g695_n_spl_
  );


  and

  (
    g697_p,
    g676_p_spl_,
    g695_n_spl_
  );


  or

  (
    g697_n,
    g676_n_spl_,
    g695_p_spl_
  );


  and

  (
    g698_p,
    g696_n_spl_,
    g697_n
  );


  or

  (
    g698_n,
    g696_p_spl_,
    g697_p
  );


  and

  (
    g699_p,
    g675_n_spl_,
    g698_p_spl_
  );


  or

  (
    g699_n,
    g675_p,
    g698_n
  );


  or

  (
    g700_n,
    g675_n_spl_,
    g698_p_spl_
  );


  and

  (
    g701_p,
    g699_n,
    g700_n
  );


  and

  (
    g702_p,
    g672_n,
    g673_p_spl_
  );


  or

  (
    g702_n,
    g672_p_spl_,
    g673_n
  );


  and

  (
    g703_p,
    n2809_lo_p_spl_000,
    n6148_o2_p_spl_0
  );


  or

  (
    g703_n,
    n2809_lo_n_spl_000,
    n6148_o2_n_spl_0
  );


  and

  (
    g704_p,
    n2734_lo_p_spl_000,
    lo002_buf_o2_p_spl_00
  );


  or

  (
    g704_n,
    n2734_lo_n_spl_000,
    lo002_buf_o2_n_spl_00
  );


  and

  (
    g705_p,
    n2045_o2_p,
    n2048_o2_n
  );


  or

  (
    g705_n,
    n2045_o2_n,
    n2048_o2_p
  );


  and

  (
    g706_p,
    n2099_o2_n_spl_,
    n2104_o2_p_spl_
  );


  or

  (
    g706_n,
    n2099_o2_p_spl_,
    n2104_o2_n_spl_
  );


  and

  (
    g707_p,
    n2099_o2_p_spl_,
    n2104_o2_n_spl_
  );


  or

  (
    g707_n,
    n2099_o2_n_spl_,
    n2104_o2_p_spl_
  );


  and

  (
    g708_p,
    g706_n_spl_,
    g707_n
  );


  or

  (
    g708_n,
    g706_p_spl_,
    g707_p
  );


  and

  (
    g709_p,
    g705_n_spl_,
    g708_p_spl_
  );


  or

  (
    g709_n,
    g705_p_spl_,
    g708_n_spl_
  );


  and

  (
    g710_p,
    n4847_o2_p_spl_0,
    lo110_buf_o2_p_spl_0
  );


  or

  (
    g710_n,
    n4847_o2_n_spl_0,
    lo110_buf_o2_n_spl_0
  );


  and

  (
    g711_p,
    g705_p_spl_,
    g708_n_spl_
  );


  or

  (
    g711_n,
    g705_n_spl_,
    g708_p_spl_
  );


  and

  (
    g712_p,
    g709_n_spl_,
    g711_n
  );


  or

  (
    g712_n,
    g709_p_spl_,
    g711_p
  );


  and

  (
    g713_p,
    g710_n_spl_,
    g712_p_spl_
  );


  or

  (
    g713_n,
    g710_p_spl_,
    g712_n_spl_
  );


  and

  (
    g714_p,
    g709_n_spl_,
    g713_n_spl_
  );


  or

  (
    g714_n,
    g709_p_spl_,
    g713_p_spl_
  );


  and

  (
    g715_p,
    n4848_o2_p_spl_0,
    lo110_buf_o2_p_spl_0
  );


  or

  (
    g715_n,
    n4848_o2_n_spl_0,
    lo110_buf_o2_n_spl_0
  );


  and

  (
    g716_p,
    n4849_o2_p_spl_0,
    lo106_buf_o2_p
  );


  or

  (
    g716_n,
    n4849_o2_n_spl_0,
    lo106_buf_o2_n
  );


  and

  (
    g717_p,
    n2102_o2_p,
    g706_n_spl_
  );


  or

  (
    g717_n,
    n2102_o2_n,
    g706_p_spl_
  );


  and

  (
    g718_p,
    g716_n_spl_,
    g717_n_spl_
  );


  or

  (
    g718_n,
    g716_p_spl_,
    g717_p_spl_
  );


  and

  (
    g719_p,
    g716_p_spl_,
    g717_p_spl_
  );


  or

  (
    g719_n,
    g716_n_spl_,
    g717_n_spl_
  );


  and

  (
    g720_p,
    g718_n_spl_,
    g719_n
  );


  or

  (
    g720_n,
    g718_p_spl_,
    g719_p
  );


  and

  (
    g721_p,
    g715_n_spl_,
    g720_p_spl_
  );


  or

  (
    g721_n,
    g715_p_spl_,
    g720_n_spl_
  );


  and

  (
    g722_p,
    g715_p_spl_,
    g720_n_spl_
  );


  or

  (
    g722_n,
    g715_n_spl_,
    g720_p_spl_
  );


  and

  (
    g723_p,
    g721_n_spl_,
    g722_n
  );


  or

  (
    g723_n,
    g721_p_spl_,
    g722_p
  );


  and

  (
    g724_p,
    g714_n_spl_,
    g723_p_spl_
  );


  or

  (
    g724_n,
    g714_p_spl_,
    g723_n_spl_
  );


  and

  (
    g725_p,
    n4847_o2_p_spl_0,
    lo114_buf_o2_p_spl_00
  );


  or

  (
    g725_n,
    n4847_o2_n_spl_0,
    lo114_buf_o2_n_spl_00
  );


  and

  (
    g726_p,
    g714_p_spl_,
    g723_n_spl_
  );


  or

  (
    g726_n,
    g714_n_spl_,
    g723_p_spl_
  );


  and

  (
    g727_p,
    g724_n_spl_,
    g726_n
  );


  or

  (
    g727_n,
    g724_p_spl_,
    g726_p
  );


  and

  (
    g728_p,
    g725_n_spl_,
    g727_p_spl_
  );


  or

  (
    g728_n,
    g725_p_spl_,
    g727_n_spl_
  );


  and

  (
    g729_p,
    g724_n_spl_,
    g728_n_spl_
  );


  or

  (
    g729_n,
    g724_p_spl_,
    g728_p_spl_
  );


  and

  (
    g730_p,
    n4848_o2_p_spl_0,
    lo114_buf_o2_p_spl_00
  );


  or

  (
    g730_n,
    n4848_o2_n_spl_0,
    lo114_buf_o2_n_spl_00
  );


  and

  (
    g731_p,
    n4849_o2_p_spl_0,
    lo110_buf_o2_p_spl_1
  );


  or

  (
    g731_n,
    n4849_o2_n_spl_0,
    lo110_buf_o2_n_spl_1
  );


  and

  (
    g732_p,
    g718_n_spl_,
    g721_n_spl_
  );


  or

  (
    g732_n,
    g718_p_spl_,
    g721_p_spl_
  );


  and

  (
    g733_p,
    g731_n_spl_,
    g732_n_spl_
  );


  or

  (
    g733_n,
    g731_p_spl_,
    g732_p_spl_
  );


  and

  (
    g734_p,
    g731_p_spl_,
    g732_p_spl_
  );


  or

  (
    g734_n,
    g731_n_spl_,
    g732_n_spl_
  );


  and

  (
    g735_p,
    g733_n_spl_,
    g734_n
  );


  or

  (
    g735_n,
    g733_p_spl_,
    g734_p
  );


  and

  (
    g736_p,
    g730_n_spl_,
    g735_p_spl_
  );


  or

  (
    g736_n,
    g730_p_spl_,
    g735_n_spl_
  );


  and

  (
    g737_p,
    g730_p_spl_,
    g735_n_spl_
  );


  or

  (
    g737_n,
    g730_n_spl_,
    g735_p_spl_
  );


  and

  (
    g738_p,
    g736_n_spl_,
    g737_n
  );


  or

  (
    g738_n,
    g736_p_spl_,
    g737_p
  );


  and

  (
    g739_p,
    g729_n_spl_,
    g738_p_spl_
  );


  or

  (
    g739_n,
    g729_p_spl_,
    g738_n_spl_
  );


  and

  (
    g740_p,
    n1913_o2_p,
    n1916_o2_n
  );


  or

  (
    g740_n,
    n1913_o2_n,
    n1916_o2_p
  );


  and

  (
    g741_p,
    n1959_o2_n_spl_,
    n1988_o2_p_spl_
  );


  or

  (
    g741_n,
    n1959_o2_p_spl_,
    n1988_o2_n_spl_
  );


  and

  (
    g742_p,
    n1959_o2_p_spl_,
    n1988_o2_n_spl_
  );


  or

  (
    g742_n,
    n1959_o2_n_spl_,
    n1988_o2_p_spl_
  );


  and

  (
    g743_p,
    g741_n_spl_,
    g742_n
  );


  or

  (
    g743_n,
    g741_p_spl_,
    g742_p
  );


  and

  (
    g744_p,
    g740_n_spl_,
    g743_p_spl_
  );


  or

  (
    g744_n,
    g740_p_spl_,
    g743_n_spl_
  );


  and

  (
    g745_p,
    n4844_o2_p_spl_0,
    lo114_buf_o2_p_spl_01
  );


  or

  (
    g745_n,
    n4844_o2_n_spl_0,
    lo114_buf_o2_n_spl_01
  );


  and

  (
    g746_p,
    g740_p_spl_,
    g743_n_spl_
  );


  or

  (
    g746_n,
    g740_n_spl_,
    g743_p_spl_
  );


  and

  (
    g747_p,
    g744_n_spl_,
    g746_n
  );


  or

  (
    g747_n,
    g744_p_spl_,
    g746_p
  );


  and

  (
    g748_p,
    g745_n_spl_,
    g747_p_spl_
  );


  or

  (
    g748_n,
    g745_p_spl_,
    g747_n_spl_
  );


  and

  (
    g749_p,
    g744_n_spl_,
    g748_n_spl_
  );


  or

  (
    g749_n,
    g744_p_spl_,
    g748_p_spl_
  );


  and

  (
    g750_p,
    n4845_o2_p_spl_0,
    lo114_buf_o2_p_spl_01
  );


  or

  (
    g750_n,
    n4845_o2_n_spl_0,
    lo114_buf_o2_n_spl_01
  );


  and

  (
    g751_p,
    n1986_o2_p,
    g741_n_spl_
  );


  or

  (
    g751_n,
    n1986_o2_n,
    g741_p_spl_
  );


  and

  (
    g752_p,
    n4846_o2_p_spl_0,
    lo110_buf_o2_p_spl_1
  );


  or

  (
    g752_n,
    n4846_o2_n_spl_0,
    lo110_buf_o2_n_spl_1
  );


  and

  (
    g753_p,
    n2033_o2_n_spl_,
    n2050_o2_n_spl_
  );


  or

  (
    g753_n,
    n2033_o2_p_spl_,
    n2050_o2_p_spl_
  );


  and

  (
    g754_p,
    n2033_o2_p_spl_,
    n2050_o2_p_spl_
  );


  or

  (
    g754_n,
    n2033_o2_n_spl_,
    n2050_o2_n_spl_
  );


  and

  (
    g755_p,
    g753_n_spl_,
    g754_n
  );


  or

  (
    g755_n,
    g753_p_spl_,
    g754_p
  );


  and

  (
    g756_p,
    g752_n_spl_,
    g755_p_spl_
  );


  or

  (
    g756_n,
    g752_p_spl_,
    g755_n_spl_
  );


  and

  (
    g757_p,
    g752_p_spl_,
    g755_n_spl_
  );


  or

  (
    g757_n,
    g752_n_spl_,
    g755_p_spl_
  );


  and

  (
    g758_p,
    g756_n_spl_,
    g757_n
  );


  or

  (
    g758_n,
    g756_p_spl_,
    g757_p
  );


  and

  (
    g759_p,
    g751_n_spl_,
    g758_p_spl_
  );


  or

  (
    g759_n,
    g751_p_spl_,
    g758_n_spl_
  );


  and

  (
    g760_p,
    g751_p_spl_,
    g758_n_spl_
  );


  or

  (
    g760_n,
    g751_n_spl_,
    g758_p_spl_
  );


  and

  (
    g761_p,
    g759_n_spl_,
    g760_n
  );


  or

  (
    g761_n,
    g759_p_spl_,
    g760_p
  );


  and

  (
    g762_p,
    g750_n_spl_,
    g761_p_spl_
  );


  or

  (
    g762_n,
    g750_p_spl_,
    g761_n_spl_
  );


  and

  (
    g763_p,
    g750_p_spl_,
    g761_n_spl_
  );


  or

  (
    g763_n,
    g750_n_spl_,
    g761_p_spl_
  );


  and

  (
    g764_p,
    g762_n_spl_,
    g763_n
  );


  or

  (
    g764_n,
    g762_p_spl_,
    g763_p
  );


  and

  (
    g765_p,
    g749_n_spl_,
    g764_p_spl_
  );


  or

  (
    g765_n,
    g749_p_spl_,
    g764_n_spl_
  );


  and

  (
    g766_p,
    n4844_o2_p_spl_0,
    lo118_buf_o2_p_spl_000
  );


  or

  (
    g766_n,
    n4844_o2_n_spl_0,
    lo118_buf_o2_n_spl_000
  );


  and

  (
    g767_p,
    g749_p_spl_,
    g764_n_spl_
  );


  or

  (
    g767_n,
    g749_n_spl_,
    g764_p_spl_
  );


  and

  (
    g768_p,
    g765_n_spl_,
    g767_n
  );


  or

  (
    g768_n,
    g765_p_spl_,
    g767_p
  );


  and

  (
    g769_p,
    g766_n_spl_,
    g768_p_spl_
  );


  or

  (
    g769_n,
    g766_p_spl_,
    g768_n_spl_
  );


  and

  (
    g770_p,
    g765_n_spl_,
    g769_n_spl_
  );


  or

  (
    g770_n,
    g765_p_spl_,
    g769_p_spl_
  );


  and

  (
    g771_p,
    n4845_o2_p_spl_0,
    lo118_buf_o2_p_spl_00
  );


  or

  (
    g771_n,
    n4845_o2_n_spl_0,
    lo118_buf_o2_n_spl_00
  );


  and

  (
    g772_p,
    g759_n_spl_,
    g762_n_spl_
  );


  or

  (
    g772_n,
    g759_p_spl_,
    g762_p_spl_
  );


  and

  (
    g773_p,
    n4846_o2_p_spl_0,
    lo114_buf_o2_p_spl_10
  );


  or

  (
    g773_n,
    n4846_o2_n_spl_0,
    lo114_buf_o2_n_spl_10
  );


  and

  (
    g774_p,
    g753_n_spl_,
    g756_n_spl_
  );


  or

  (
    g774_n,
    g753_p_spl_,
    g756_p_spl_
  );


  and

  (
    g775_p,
    g710_p_spl_,
    g712_n_spl_
  );


  or

  (
    g775_n,
    g710_n_spl_,
    g712_p_spl_
  );


  and

  (
    g776_p,
    g713_n_spl_,
    g775_n
  );


  or

  (
    g776_n,
    g713_p_spl_,
    g775_p
  );


  and

  (
    g777_p,
    g774_n_spl_,
    g776_p_spl_
  );


  or

  (
    g777_n,
    g774_p_spl_,
    g776_n_spl_
  );


  and

  (
    g778_p,
    g774_p_spl_,
    g776_n_spl_
  );


  or

  (
    g778_n,
    g774_n_spl_,
    g776_p_spl_
  );


  and

  (
    g779_p,
    g777_n_spl_,
    g778_n
  );


  or

  (
    g779_n,
    g777_p_spl_,
    g778_p
  );


  and

  (
    g780_p,
    g773_n_spl_,
    g779_p_spl_
  );


  or

  (
    g780_n,
    g773_p_spl_,
    g779_n_spl_
  );


  and

  (
    g781_p,
    g773_p_spl_,
    g779_n_spl_
  );


  or

  (
    g781_n,
    g773_n_spl_,
    g779_p_spl_
  );


  and

  (
    g782_p,
    g780_n_spl_,
    g781_n
  );


  or

  (
    g782_n,
    g780_p_spl_,
    g781_p
  );


  and

  (
    g783_p,
    g772_n_spl_,
    g782_p_spl_
  );


  or

  (
    g783_n,
    g772_p_spl_,
    g782_n_spl_
  );


  and

  (
    g784_p,
    g772_p_spl_,
    g782_n_spl_
  );


  or

  (
    g784_n,
    g772_n_spl_,
    g782_p_spl_
  );


  and

  (
    g785_p,
    g783_n_spl_,
    g784_n
  );


  or

  (
    g785_n,
    g783_p_spl_,
    g784_p
  );


  and

  (
    g786_p,
    g771_n_spl_,
    g785_p_spl_
  );


  or

  (
    g786_n,
    g771_p_spl_,
    g785_n_spl_
  );


  and

  (
    g787_p,
    g771_p_spl_,
    g785_n_spl_
  );


  or

  (
    g787_n,
    g771_n_spl_,
    g785_p_spl_
  );


  and

  (
    g788_p,
    g786_n_spl_,
    g787_n
  );


  or

  (
    g788_n,
    g786_p_spl_,
    g787_p
  );


  and

  (
    g789_p,
    g770_n_spl_,
    g788_p_spl_
  );


  or

  (
    g789_n,
    g770_p_spl_,
    g788_n_spl_
  );


  and

  (
    g790_p,
    n1749_o2_p,
    n1752_o2_n
  );


  or

  (
    g790_n,
    n1749_o2_n,
    n1752_o2_p
  );


  and

  (
    g791_p,
    n1787_o2_n_spl_,
    n1840_o2_p_spl_
  );


  or

  (
    g791_n,
    n1787_o2_p_spl_,
    n1840_o2_n_spl_
  );


  and

  (
    g792_p,
    n1787_o2_p_spl_,
    n1840_o2_n_spl_
  );


  or

  (
    g792_n,
    n1787_o2_n_spl_,
    n1840_o2_p_spl_
  );


  and

  (
    g793_p,
    g791_n_spl_,
    g792_n
  );


  or

  (
    g793_n,
    g791_p_spl_,
    g792_p
  );


  and

  (
    g794_p,
    g790_n_spl_,
    g793_p_spl_
  );


  or

  (
    g794_n,
    g790_p_spl_,
    g793_n_spl_
  );


  and

  (
    g795_p,
    n4841_o2_p_spl_0,
    lo118_buf_o2_p_spl_01
  );


  or

  (
    g795_n,
    n4841_o2_n_spl_0,
    lo118_buf_o2_n_spl_01
  );


  and

  (
    g796_p,
    g790_p_spl_,
    g793_n_spl_
  );


  or

  (
    g796_n,
    g790_n_spl_,
    g793_p_spl_
  );


  and

  (
    g797_p,
    g794_n_spl_,
    g796_n
  );


  or

  (
    g797_n,
    g794_p_spl_,
    g796_p
  );


  and

  (
    g798_p,
    g795_n_spl_,
    g797_p_spl_
  );


  or

  (
    g798_n,
    g795_p_spl_,
    g797_n_spl_
  );


  and

  (
    g799_p,
    g794_n_spl_,
    g798_n_spl_
  );


  or

  (
    g799_n,
    g794_p_spl_,
    g798_p_spl_
  );


  and

  (
    g800_p,
    n4842_o2_p_spl_,
    lo118_buf_o2_p_spl_01
  );


  or

  (
    g800_n,
    n4842_o2_n_spl_0,
    lo118_buf_o2_n_spl_01
  );


  and

  (
    g801_p,
    n1838_o2_p,
    g791_n_spl_
  );


  or

  (
    g801_n,
    n1838_o2_n,
    g791_p_spl_
  );


  and

  (
    g802_p,
    n4843_o2_p_spl_0,
    lo114_buf_o2_p_spl_10
  );


  or

  (
    g802_n,
    n4843_o2_n_spl_0,
    lo114_buf_o2_n_spl_10
  );


  and

  (
    g803_p,
    n1877_o2_n_spl_,
    n1918_o2_n_spl_
  );


  or

  (
    g803_n,
    n1877_o2_p_spl_,
    n1918_o2_p_spl_
  );


  and

  (
    g804_p,
    n1877_o2_p_spl_,
    n1918_o2_p_spl_
  );


  or

  (
    g804_n,
    n1877_o2_n_spl_,
    n1918_o2_n_spl_
  );


  and

  (
    g805_p,
    g803_n_spl_,
    g804_n
  );


  or

  (
    g805_n,
    g803_p_spl_,
    g804_p
  );


  and

  (
    g806_p,
    g802_n_spl_,
    g805_p_spl_
  );


  or

  (
    g806_n,
    g802_p_spl_,
    g805_n_spl_
  );


  and

  (
    g807_p,
    g802_p_spl_,
    g805_n_spl_
  );


  or

  (
    g807_n,
    g802_n_spl_,
    g805_p_spl_
  );


  and

  (
    g808_p,
    g806_n_spl_,
    g807_n
  );


  or

  (
    g808_n,
    g806_p_spl_,
    g807_p
  );


  and

  (
    g809_p,
    g801_n_spl_,
    g808_p_spl_
  );


  or

  (
    g809_n,
    g801_p_spl_,
    g808_n_spl_
  );


  and

  (
    g810_p,
    g801_p_spl_,
    g808_n_spl_
  );


  or

  (
    g810_n,
    g801_n_spl_,
    g808_p_spl_
  );


  and

  (
    g811_p,
    g809_n_spl_,
    g810_n
  );


  or

  (
    g811_n,
    g809_p_spl_,
    g810_p
  );


  and

  (
    g812_p,
    g800_n_spl_,
    g811_p_spl_
  );


  or

  (
    g812_n,
    g800_p_spl_,
    g811_n_spl_
  );


  and

  (
    g813_p,
    g800_p_spl_,
    g811_n_spl_
  );


  or

  (
    g813_n,
    g800_n_spl_,
    g811_p_spl_
  );


  and

  (
    g814_p,
    g812_n_spl_,
    g813_n
  );


  or

  (
    g814_n,
    g812_p_spl_,
    g813_p
  );


  and

  (
    g815_p,
    g799_n_spl_,
    g814_p_spl_
  );


  or

  (
    g815_n,
    g799_p_spl_,
    g814_n_spl_
  );


  and

  (
    g816_p,
    n2848_lo_p_spl_011,
    n4841_o2_p_spl_0
  );


  or

  (
    g816_n,
    n2848_lo_n_spl_011,
    n4841_o2_n_spl_0
  );


  and

  (
    g817_p,
    g799_p_spl_,
    g814_n_spl_
  );


  or

  (
    g817_n,
    g799_n_spl_,
    g814_p_spl_
  );


  and

  (
    g818_p,
    g815_n_spl_,
    g817_n
  );


  or

  (
    g818_n,
    g815_p_spl_,
    g817_p
  );


  and

  (
    g819_p,
    g816_n_spl_,
    g818_p_spl_
  );


  or

  (
    g819_n,
    g816_p_spl_,
    g818_n_spl_
  );


  and

  (
    g820_p,
    g815_n_spl_,
    g819_n_spl_
  );


  or

  (
    g820_n,
    g815_p_spl_,
    g819_p_spl_
  );


  and

  (
    g821_p,
    n2848_lo_p_spl_011,
    n4842_o2_p_spl_
  );


  or

  (
    g821_n,
    n2848_lo_n_spl_011,
    n4842_o2_n_spl_0
  );


  and

  (
    g822_p,
    g809_n_spl_,
    g812_n_spl_
  );


  or

  (
    g822_n,
    g809_p_spl_,
    g812_p_spl_
  );


  and

  (
    g823_p,
    n4843_o2_p_spl_0,
    lo118_buf_o2_p_spl_10
  );


  or

  (
    g823_n,
    n4843_o2_n_spl_0,
    lo118_buf_o2_n_spl_10
  );


  and

  (
    g824_p,
    g803_n_spl_,
    g806_n_spl_
  );


  or

  (
    g824_n,
    g803_p_spl_,
    g806_p_spl_
  );


  and

  (
    g825_p,
    g745_p_spl_,
    g747_n_spl_
  );


  or

  (
    g825_n,
    g745_n_spl_,
    g747_p_spl_
  );


  and

  (
    g826_p,
    g748_n_spl_,
    g825_n
  );


  or

  (
    g826_n,
    g748_p_spl_,
    g825_p
  );


  and

  (
    g827_p,
    g824_n_spl_,
    g826_p_spl_
  );


  or

  (
    g827_n,
    g824_p_spl_,
    g826_n_spl_
  );


  and

  (
    g828_p,
    g824_p_spl_,
    g826_n_spl_
  );


  or

  (
    g828_n,
    g824_n_spl_,
    g826_p_spl_
  );


  and

  (
    g829_p,
    g827_n_spl_,
    g828_n
  );


  or

  (
    g829_n,
    g827_p_spl_,
    g828_p
  );


  and

  (
    g830_p,
    g823_n_spl_,
    g829_p_spl_
  );


  or

  (
    g830_n,
    g823_p_spl_,
    g829_n_spl_
  );


  and

  (
    g831_p,
    g823_p_spl_,
    g829_n_spl_
  );


  or

  (
    g831_n,
    g823_n_spl_,
    g829_p_spl_
  );


  and

  (
    g832_p,
    g830_n_spl_,
    g831_n
  );


  or

  (
    g832_n,
    g830_p_spl_,
    g831_p
  );


  and

  (
    g833_p,
    g822_n_spl_,
    g832_p_spl_
  );


  or

  (
    g833_n,
    g822_p_spl_,
    g832_n_spl_
  );


  and

  (
    g834_p,
    g822_p_spl_,
    g832_n_spl_
  );


  or

  (
    g834_n,
    g822_n_spl_,
    g832_p_spl_
  );


  and

  (
    g835_p,
    g833_n_spl_,
    g834_n
  );


  or

  (
    g835_n,
    g833_p_spl_,
    g834_p
  );


  and

  (
    g836_p,
    g821_n_spl_,
    g835_p_spl_
  );


  or

  (
    g836_n,
    g821_p_spl_,
    g835_n_spl_
  );


  and

  (
    g837_p,
    g821_p_spl_,
    g835_n_spl_
  );


  or

  (
    g837_n,
    g821_n_spl_,
    g835_p_spl_
  );


  and

  (
    g838_p,
    g836_n_spl_,
    g837_n
  );


  or

  (
    g838_n,
    g836_p_spl_,
    g837_p
  );


  and

  (
    g839_p,
    g820_n_spl_,
    g838_p_spl_
  );


  or

  (
    g839_n,
    g820_p_spl_,
    g838_n_spl_
  );


  and

  (
    g840_p,
    g674_n_spl_,
    g701_p_spl_
  );


  and

  (
    g841_p,
    g668_n_spl_,
    g671_n
  );


  or

  (
    g841_n,
    g668_p_spl_,
    g671_p_spl_
  );


  and

  (
    g842_p,
    n2797_lo_p_spl_000,
    n6053_o2_p_spl_00
  );


  or

  (
    g842_n,
    n2797_lo_n_spl_000,
    n6053_o2_n_spl_00
  );


  and

  (
    g843_p,
    n839_o2_p_spl_,
    g665_n_spl_
  );


  or

  (
    g843_n,
    n839_o2_n_spl_,
    g665_p_spl_
  );


  and

  (
    g844_p,
    n6024_o2_p_spl_00,
    lo102_buf_o2_p_spl_001
  );


  or

  (
    g844_n,
    n6024_o2_n_spl_00,
    lo102_buf_o2_n_spl_001
  );


  and

  (
    g845_p,
    n917_o2_p_spl_,
    n918_o2_n
  );


  or

  (
    g845_n,
    n917_o2_n_spl_,
    n918_o2_p
  );


  and

  (
    g846_p,
    g844_n_spl_,
    g845_p_spl_
  );


  or

  (
    g846_n,
    g844_p_spl_,
    g845_n_spl_
  );


  and

  (
    g847_p,
    g844_p_spl_,
    g845_n_spl_
  );


  or

  (
    g847_n,
    g844_n_spl_,
    g845_p_spl_
  );


  and

  (
    g848_p,
    g846_n_spl_,
    g847_n
  );


  or

  (
    g848_n,
    g846_p_spl_,
    g847_p
  );


  and

  (
    g849_p,
    g843_n_spl_,
    g848_p_spl_
  );


  or

  (
    g849_n,
    g843_p_spl_,
    g848_n_spl_
  );


  and

  (
    g850_p,
    g843_p_spl_,
    g848_n_spl_
  );


  or

  (
    g850_n,
    g843_n_spl_,
    g848_p_spl_
  );


  and

  (
    g851_p,
    g849_n_spl_,
    g850_n
  );


  or

  (
    g851_n,
    g849_p_spl_,
    g850_p
  );


  and

  (
    g852_p,
    g842_n_spl_,
    g851_p_spl_
  );


  or

  (
    g852_n,
    g842_p_spl_,
    g851_n_spl_
  );


  and

  (
    g853_p,
    g842_p_spl_,
    g851_n_spl_
  );


  or

  (
    g853_n,
    g842_n_spl_,
    g851_p_spl_
  );


  and

  (
    g854_p,
    g852_n_spl_,
    g853_n
  );


  or

  (
    g854_n,
    g852_p_spl_,
    g853_p
  );


  and

  (
    g855_p,
    g841_n_spl_,
    g854_p_spl_
  );


  or

  (
    g855_n,
    g841_p_spl_,
    g854_n_spl_
  );


  and

  (
    g856_p,
    g841_p_spl_,
    g854_n_spl_
  );


  or

  (
    g856_n,
    g841_n_spl_,
    g854_p_spl_
  );


  and

  (
    g857_p,
    g855_n_spl_,
    g856_n
  );


  or

  (
    g857_n,
    g855_p_spl_,
    g856_p
  );


  and

  (
    g858_p,
    n509_o2_p_spl_,
    g702_n
  );


  or

  (
    g858_n,
    n509_o2_n_spl_,
    g702_p_spl_
  );


  and

  (
    g859_p,
    n517_o2_n_spl_,
    n541_o2_p_spl_
  );


  or

  (
    g859_n,
    n517_o2_p_spl_,
    n541_o2_n_spl_
  );


  and

  (
    g860_p,
    n517_o2_p_spl_,
    n541_o2_n_spl_
  );


  or

  (
    g860_n,
    n517_o2_n_spl_,
    n541_o2_p_spl_
  );


  and

  (
    g861_p,
    g859_n_spl_,
    g860_n
  );


  or

  (
    g861_n,
    g859_p_spl_,
    g860_p
  );


  and

  (
    g862_p,
    g858_n_spl_,
    g861_p_spl_
  );


  or

  (
    g862_n,
    g858_p_spl_,
    g861_n_spl_
  );


  and

  (
    g863_p,
    g858_p_spl_,
    g861_n_spl_
  );


  or

  (
    g863_n,
    g858_n_spl_,
    g861_p_spl_
  );


  and

  (
    g864_p,
    g862_n_spl_,
    g863_n
  );


  or

  (
    g864_n,
    g862_p_spl_,
    g863_p
  );


  and

  (
    g865_p,
    g703_n,
    g857_p_spl_
  );


  or

  (
    g865_n,
    g703_p_spl_,
    g857_n
  );


  and

  (
    g866_p,
    g704_n,
    g864_p_spl_
  );


  or

  (
    g866_n,
    g704_p_spl_,
    g864_n
  );


  or

  (
    g867_n,
    g699_p,
    g840_p_spl_
  );


  and

  (
    g868_p,
    g693_n_spl_,
    g696_n_spl_
  );


  or

  (
    g868_n,
    g693_p_spl_,
    g696_p_spl_
  );


  and

  (
    g869_p,
    n2860_lo_p_spl_10,
    n4839_o2_p_spl_
  );


  or

  (
    g869_n,
    n2860_lo_n_spl_10,
    n4839_o2_n_spl_
  );


  and

  (
    g870_p,
    g687_n_spl_,
    g690_n_spl_
  );


  or

  (
    g870_n,
    g687_p_spl_,
    g690_p_spl_
  );


  and

  (
    g871_p,
    n2848_lo_p_spl_10,
    n4840_o2_p_spl_0
  );


  or

  (
    g871_n,
    n2848_lo_n_spl_10,
    n4840_o2_n_spl_0
  );


  and

  (
    g872_p,
    g681_n_spl_,
    g684_n_spl_
  );


  or

  (
    g872_n,
    g681_p_spl_,
    g684_p_spl_
  );


  and

  (
    g873_p,
    g795_p_spl_,
    g797_n_spl_
  );


  or

  (
    g873_n,
    g795_n_spl_,
    g797_p_spl_
  );


  and

  (
    g874_p,
    g798_n_spl_,
    g873_n
  );


  or

  (
    g874_n,
    g798_p_spl_,
    g873_p
  );


  and

  (
    g875_p,
    g872_n_spl_,
    g874_p_spl_
  );


  or

  (
    g875_n,
    g872_p_spl_,
    g874_n_spl_
  );


  and

  (
    g876_p,
    g872_p_spl_,
    g874_n_spl_
  );


  or

  (
    g876_n,
    g872_n_spl_,
    g874_p_spl_
  );


  and

  (
    g877_p,
    g875_n_spl_,
    g876_n
  );


  or

  (
    g877_n,
    g875_p_spl_,
    g876_p
  );


  and

  (
    g878_p,
    g871_n_spl_,
    g877_p_spl_
  );


  or

  (
    g878_n,
    g871_p_spl_,
    g877_n_spl_
  );


  and

  (
    g879_p,
    g871_p_spl_,
    g877_n_spl_
  );


  or

  (
    g879_n,
    g871_n_spl_,
    g877_p_spl_
  );


  and

  (
    g880_p,
    g878_n_spl_,
    g879_n
  );


  or

  (
    g880_n,
    g878_p_spl_,
    g879_p
  );


  and

  (
    g881_p,
    g870_n_spl_,
    g880_p_spl_
  );


  or

  (
    g881_n,
    g870_p_spl_,
    g880_n_spl_
  );


  and

  (
    g882_p,
    g870_p_spl_,
    g880_n_spl_
  );


  or

  (
    g882_n,
    g870_n_spl_,
    g880_p_spl_
  );


  and

  (
    g883_p,
    g881_n_spl_,
    g882_n
  );


  or

  (
    g883_n,
    g881_p_spl_,
    g882_p
  );


  and

  (
    g884_p,
    g869_n_spl_,
    g883_p_spl_
  );


  or

  (
    g884_n,
    g869_p_spl_,
    g883_n_spl_
  );


  and

  (
    g885_p,
    g869_p_spl_,
    g883_n_spl_
  );


  or

  (
    g885_n,
    g869_n_spl_,
    g883_p_spl_
  );


  and

  (
    g886_p,
    g884_n_spl_,
    g885_n
  );


  or

  (
    g886_n,
    g884_p_spl_,
    g885_p
  );


  and

  (
    g887_p,
    g868_n_spl_,
    g886_p_spl_
  );


  or

  (
    g887_n,
    g868_p,
    g886_n
  );


  or

  (
    g888_n,
    g868_n_spl_,
    g886_p_spl_
  );


  and

  (
    g889_p,
    g887_n,
    g888_n
  );


  and

  (
    g890_p,
    n2746_lo_p_spl_000,
    lo002_buf_o2_p_spl_0
  );


  or

  (
    g890_n,
    n2746_lo_n_spl_000,
    lo002_buf_o2_n_spl_0
  );


  and

  (
    g891_p,
    g862_n_spl_,
    g866_n
  );


  or

  (
    g891_n,
    g862_p_spl_,
    g866_p_spl_
  );


  and

  (
    g892_p,
    n2734_lo_p_spl_000,
    lo006_buf_o2_p_spl_00
  );


  or

  (
    g892_n,
    n2734_lo_n_spl_000,
    lo006_buf_o2_n_spl_0
  );


  and

  (
    g893_p,
    n539_o2_p,
    g859_n_spl_
  );


  or

  (
    g893_n,
    n539_o2_n,
    g859_p_spl_
  );


  and

  (
    g894_p,
    n555_o2_n_spl_,
    n579_o2_p_spl_
  );


  or

  (
    g894_n,
    n555_o2_p_spl_,
    n579_o2_n_spl_
  );


  and

  (
    g895_p,
    n555_o2_p_spl_,
    n579_o2_n_spl_
  );


  or

  (
    g895_n,
    n555_o2_n_spl_,
    n579_o2_p_spl_
  );


  and

  (
    g896_p,
    g894_n_spl_,
    g895_n
  );


  or

  (
    g896_n,
    g894_p_spl_,
    g895_p
  );


  and

  (
    g897_p,
    g893_n_spl_,
    g896_p_spl_
  );


  or

  (
    g897_n,
    g893_p_spl_,
    g896_n_spl_
  );


  and

  (
    g898_p,
    g893_p_spl_,
    g896_n_spl_
  );


  or

  (
    g898_n,
    g893_n_spl_,
    g896_p_spl_
  );


  and

  (
    g899_p,
    g897_n_spl_,
    g898_n
  );


  or

  (
    g899_n,
    g897_p_spl_,
    g898_p
  );


  and

  (
    g900_p,
    g892_n_spl_,
    g899_p_spl_
  );


  or

  (
    g900_n,
    g892_p_spl_,
    g899_n_spl_
  );


  and

  (
    g901_p,
    g892_p_spl_,
    g899_n_spl_
  );


  or

  (
    g901_n,
    g892_n_spl_,
    g899_p_spl_
  );


  and

  (
    g902_p,
    g900_n_spl_,
    g901_n
  );


  or

  (
    g902_n,
    g900_p_spl_,
    g901_p
  );


  and

  (
    g903_p,
    g891_n_spl_,
    g902_p_spl_
  );


  or

  (
    g903_n,
    g891_p_spl_,
    g902_n_spl_
  );


  and

  (
    g904_p,
    g891_p_spl_,
    g902_n_spl_
  );


  or

  (
    g904_n,
    g891_n_spl_,
    g902_p_spl_
  );


  and

  (
    g905_p,
    g903_n_spl_,
    g904_n
  );


  or

  (
    g905_n,
    g903_p_spl_,
    g904_p
  );


  and

  (
    g906_p,
    g890_n,
    g905_p_spl_
  );


  or

  (
    g906_n,
    g890_p_spl_,
    g905_n
  );


  and

  (
    g907_p,
    n2821_lo_p_spl_000,
    n6148_o2_p_spl_1
  );


  or

  (
    g907_n,
    n2821_lo_n_spl_00,
    n6148_o2_n_spl_1
  );


  and

  (
    g908_p,
    n2860_lo_p_spl_10,
    n4841_o2_p_spl_
  );


  or

  (
    g908_n,
    n2860_lo_n_spl_10,
    n4841_o2_n_spl_
  );


  and

  (
    g909_p,
    g820_p_spl_,
    g838_n_spl_
  );


  or

  (
    g909_n,
    g820_n_spl_,
    g838_p_spl_
  );


  and

  (
    g910_p,
    g839_n_spl_,
    g909_n
  );


  or

  (
    g910_n,
    g839_p,
    g909_p
  );


  or

  (
    g911_n,
    g908_p,
    g910_n
  );


  and

  (
    g912_p,
    n2848_lo_p_spl_10,
    n4844_o2_p_spl_1
  );


  or

  (
    g912_n,
    n2848_lo_n_spl_10,
    n4844_o2_n_spl_
  );


  and

  (
    g913_p,
    g770_p_spl_,
    g788_n_spl_
  );


  or

  (
    g913_n,
    g770_n_spl_,
    g788_p_spl_
  );


  and

  (
    g914_p,
    g789_n_spl_,
    g913_n
  );


  or

  (
    g914_n,
    g789_p,
    g913_p
  );


  or

  (
    g915_n,
    g912_p,
    g914_n
  );


  and

  (
    g916_p,
    n4847_o2_p_spl_1,
    lo118_buf_o2_p_spl_10
  );


  or

  (
    g916_n,
    n4847_o2_n_spl_,
    lo118_buf_o2_n_spl_10
  );


  and

  (
    g917_p,
    g729_p_spl_,
    g738_n_spl_
  );


  or

  (
    g917_n,
    g729_n_spl_,
    g738_p_spl_
  );


  and

  (
    g918_p,
    g739_n_spl_,
    g917_n
  );


  or

  (
    g918_n,
    g739_p,
    g917_p
  );


  or

  (
    g919_n,
    g916_p,
    g918_n
  );


  and

  (
    g920_p,
    n4849_o2_p_spl_1,
    lo114_buf_o2_p_spl_1
  );


  or

  (
    g920_n,
    n4849_o2_n_spl_,
    lo114_buf_o2_n_spl_1
  );


  and

  (
    g921_p,
    g733_n_spl_,
    g736_n_spl_
  );


  or

  (
    g921_n,
    g733_p_spl_,
    g736_p_spl_
  );


  or

  (
    g922_n,
    g920_p,
    g921_p
  );


  and

  (
    g923_p,
    g783_n_spl_,
    g786_n_spl_
  );


  or

  (
    g923_n,
    g783_p_spl_,
    g786_p_spl_
  );


  and

  (
    g924_p,
    n4846_o2_p_spl_1,
    lo118_buf_o2_p_spl_11
  );


  or

  (
    g924_n,
    n4846_o2_n_spl_,
    lo118_buf_o2_n_spl_11
  );


  and

  (
    g925_p,
    g777_n_spl_,
    g780_n_spl_
  );


  or

  (
    g925_n,
    g777_p_spl_,
    g780_p_spl_
  );


  and

  (
    g926_p,
    g725_p_spl_,
    g727_n_spl_
  );


  or

  (
    g926_n,
    g725_n_spl_,
    g727_p_spl_
  );


  and

  (
    g927_p,
    g728_n_spl_,
    g926_n
  );


  or

  (
    g927_n,
    g728_p_spl_,
    g926_p
  );


  and

  (
    g928_p,
    g925_n_spl_,
    g927_p_spl_
  );


  or

  (
    g928_n,
    g925_p_spl_,
    g927_n_spl_
  );


  and

  (
    g929_p,
    g925_p_spl_,
    g927_n_spl_
  );


  or

  (
    g929_n,
    g925_n_spl_,
    g927_p_spl_
  );


  and

  (
    g930_p,
    g928_n,
    g929_n
  );


  or

  (
    g930_n,
    g928_p_spl_,
    g929_p
  );


  and

  (
    g931_p,
    g924_n_spl_,
    g930_p_spl_
  );


  or

  (
    g931_n,
    g924_p_spl_,
    g930_n_spl_
  );


  and

  (
    g932_p,
    g924_p_spl_,
    g930_n_spl_
  );


  or

  (
    g932_n,
    g924_n_spl_,
    g930_p_spl_
  );


  and

  (
    g933_p,
    g931_n,
    g932_n
  );


  or

  (
    g933_n,
    g931_p_spl_,
    g932_p
  );


  or

  (
    g934_n,
    g923_p,
    g933_n
  );


  and

  (
    g935_p,
    g833_n_spl_,
    g836_n_spl_
  );


  or

  (
    g935_n,
    g833_p_spl_,
    g836_p_spl_
  );


  and

  (
    g936_p,
    n2848_lo_p_spl_11,
    n4843_o2_p_spl_1
  );


  or

  (
    g936_n,
    n2848_lo_n_spl_11,
    n4843_o2_n_spl_
  );


  and

  (
    g937_p,
    g827_n_spl_,
    g830_n_spl_
  );


  or

  (
    g937_n,
    g827_p_spl_,
    g830_p_spl_
  );


  and

  (
    g938_p,
    g766_p_spl_,
    g768_n_spl_
  );


  or

  (
    g938_n,
    g766_n_spl_,
    g768_p_spl_
  );


  and

  (
    g939_p,
    g769_n_spl_,
    g938_n
  );


  or

  (
    g939_n,
    g769_p_spl_,
    g938_p
  );


  and

  (
    g940_p,
    g937_n_spl_,
    g939_p_spl_
  );


  or

  (
    g940_n,
    g937_p_spl_,
    g939_n_spl_
  );


  and

  (
    g941_p,
    g937_p_spl_,
    g939_n_spl_
  );


  or

  (
    g941_n,
    g937_n_spl_,
    g939_p_spl_
  );


  and

  (
    g942_p,
    g940_n,
    g941_n
  );


  or

  (
    g942_n,
    g940_p_spl_,
    g941_p
  );


  and

  (
    g943_p,
    g936_n_spl_,
    g942_p_spl_
  );


  or

  (
    g943_n,
    g936_p_spl_,
    g942_n_spl_
  );


  and

  (
    g944_p,
    g936_p_spl_,
    g942_n_spl_
  );


  or

  (
    g944_n,
    g936_n_spl_,
    g942_p_spl_
  );


  and

  (
    g945_p,
    g943_n,
    g944_n
  );


  or

  (
    g945_n,
    g943_p_spl_,
    g944_p
  );


  or

  (
    g946_n,
    g935_p,
    g945_n
  );


  and

  (
    g947_p,
    g881_n_spl_,
    g884_n_spl_
  );


  or

  (
    g947_n,
    g881_p_spl_,
    g884_p_spl_
  );


  and

  (
    g948_p,
    n2860_lo_p_spl_11,
    n4840_o2_p_spl_
  );


  or

  (
    g948_n,
    n2860_lo_n_spl_11,
    n4840_o2_n_spl_
  );


  and

  (
    g949_p,
    g875_n_spl_,
    g878_n_spl_
  );


  or

  (
    g949_n,
    g875_p_spl_,
    g878_p_spl_
  );


  and

  (
    g950_p,
    g816_p_spl_,
    g818_n_spl_
  );


  or

  (
    g950_n,
    g816_n_spl_,
    g818_p_spl_
  );


  and

  (
    g951_p,
    g819_n_spl_,
    g950_n
  );


  or

  (
    g951_n,
    g819_p_spl_,
    g950_p
  );


  and

  (
    g952_p,
    g949_n_spl_,
    g951_p_spl_
  );


  or

  (
    g952_n,
    g949_p_spl_,
    g951_n_spl_
  );


  and

  (
    g953_p,
    g949_p_spl_,
    g951_n_spl_
  );


  or

  (
    g953_n,
    g949_n_spl_,
    g951_p_spl_
  );


  and

  (
    g954_p,
    g952_n,
    g953_n
  );


  or

  (
    g954_n,
    g952_p_spl_,
    g953_p
  );


  and

  (
    g955_p,
    g948_n_spl_,
    g954_p_spl_
  );


  or

  (
    g955_n,
    g948_p_spl_,
    g954_n_spl_
  );


  and

  (
    g956_p,
    g948_p_spl_,
    g954_n_spl_
  );


  or

  (
    g956_n,
    g948_n_spl_,
    g954_p_spl_
  );


  and

  (
    g957_p,
    g955_n,
    g956_n
  );


  or

  (
    g957_n,
    g955_p_spl_,
    g956_p
  );


  or

  (
    g958_n,
    g947_p,
    g957_n
  );


  and

  (
    g959_p,
    g867_n_spl_,
    g889_p_spl_
  );


  and

  (
    g960_p,
    g855_n_spl_,
    g865_n
  );


  or

  (
    g960_n,
    g855_p_spl_,
    g865_p_spl_
  );


  and

  (
    g961_p,
    n2809_lo_p_spl_000,
    n6053_o2_p_spl_0
  );


  or

  (
    g961_n,
    n2809_lo_n_spl_000,
    n6053_o2_n_spl_0
  );


  and

  (
    g962_p,
    g849_n_spl_,
    g852_n_spl_
  );


  or

  (
    g962_n,
    g849_p_spl_,
    g852_p_spl_
  );


  and

  (
    g963_p,
    n2797_lo_p_spl_001,
    n6024_o2_p_spl_00
  );


  or

  (
    g963_n,
    n2797_lo_n_spl_001,
    n6024_o2_n_spl_00
  );


  and

  (
    g964_p,
    n917_o2_p_spl_,
    g846_n_spl_
  );


  or

  (
    g964_n,
    n917_o2_n_spl_,
    g846_p_spl_
  );


  and

  (
    g965_p,
    n6025_o2_p_spl_00,
    lo102_buf_o2_p_spl_001
  );


  or

  (
    g965_n,
    n6025_o2_n_spl_00,
    lo102_buf_o2_n_spl_001
  );


  and

  (
    g966_p,
    n1003_o2_p_spl_,
    n1004_o2_n
  );


  or

  (
    g966_n,
    n1003_o2_n_spl_,
    n1004_o2_p
  );


  and

  (
    g967_p,
    g965_n_spl_,
    g966_p_spl_
  );


  or

  (
    g967_n,
    g965_p_spl_,
    g966_n_spl_
  );


  and

  (
    g968_p,
    g965_p_spl_,
    g966_n_spl_
  );


  or

  (
    g968_n,
    g965_n_spl_,
    g966_p_spl_
  );


  and

  (
    g969_p,
    g967_n_spl_,
    g968_n
  );


  or

  (
    g969_n,
    g967_p_spl_,
    g968_p
  );


  and

  (
    g970_p,
    g964_n_spl_,
    g969_p_spl_
  );


  or

  (
    g970_n,
    g964_p_spl_,
    g969_n_spl_
  );


  and

  (
    g971_p,
    g964_p_spl_,
    g969_n_spl_
  );


  or

  (
    g971_n,
    g964_n_spl_,
    g969_p_spl_
  );


  and

  (
    g972_p,
    g970_n_spl_,
    g971_n
  );


  or

  (
    g972_n,
    g970_p_spl_,
    g971_p
  );


  and

  (
    g973_p,
    g963_n_spl_,
    g972_p_spl_
  );


  or

  (
    g973_n,
    g963_p_spl_,
    g972_n_spl_
  );


  and

  (
    g974_p,
    g963_p_spl_,
    g972_n_spl_
  );


  or

  (
    g974_n,
    g963_n_spl_,
    g972_p_spl_
  );


  and

  (
    g975_p,
    g973_n_spl_,
    g974_n
  );


  or

  (
    g975_n,
    g973_p_spl_,
    g974_p
  );


  and

  (
    g976_p,
    g962_n_spl_,
    g975_p_spl_
  );


  or

  (
    g976_n,
    g962_p_spl_,
    g975_n_spl_
  );


  and

  (
    g977_p,
    g962_p_spl_,
    g975_n_spl_
  );


  or

  (
    g977_n,
    g962_n_spl_,
    g975_p_spl_
  );


  and

  (
    g978_p,
    g976_n_spl_,
    g977_n
  );


  or

  (
    g978_n,
    g976_p_spl_,
    g977_p
  );


  and

  (
    g979_p,
    g961_n_spl_,
    g978_p_spl_
  );


  or

  (
    g979_n,
    g961_p_spl_,
    g978_n_spl_
  );


  and

  (
    g980_p,
    g961_p_spl_,
    g978_n_spl_
  );


  or

  (
    g980_n,
    g961_n_spl_,
    g978_p_spl_
  );


  and

  (
    g981_p,
    g979_n_spl_,
    g980_n
  );


  or

  (
    g981_n,
    g979_p_spl_,
    g980_p
  );


  and

  (
    g982_p,
    g960_n_spl_,
    g981_p_spl_
  );


  or

  (
    g982_n,
    g960_p_spl_,
    g981_n_spl_
  );


  and

  (
    g983_p,
    g960_p_spl_,
    g981_n_spl_
  );


  or

  (
    g983_n,
    g960_n_spl_,
    g981_p_spl_
  );


  and

  (
    g984_p,
    g982_n_spl_,
    g983_n
  );


  or

  (
    g984_n,
    g982_p_spl_,
    g983_p
  );


  and

  (
    g985_p,
    G2_p_spl_00,
    G17_p_spl_000
  );


  or

  (
    g985_n,
    G2_n_spl_0,
    G17_n_spl_000
  );


  and

  (
    g986_p,
    G1_p_spl_0,
    G18_p_spl_000
  );


  or

  (
    g986_n,
    G1_n_spl_0,
    G18_n_spl_000
  );


  and

  (
    g987_p,
    g907_n,
    g984_p_spl_
  );


  or

  (
    g987_n,
    g907_p_spl_,
    g984_n
  );


  and

  (
    g988_p,
    n2758_lo_p_spl_000,
    lo002_buf_o2_p_spl_1
  );


  or

  (
    g988_n,
    n2758_lo_n_spl_000,
    lo002_buf_o2_n_spl_1
  );


  and

  (
    g989_p,
    g985_p_spl_,
    g986_p_spl_
  );


  or

  (
    g989_n,
    g985_n,
    g986_n
  );


  and

  (
    g990_p,
    g903_n_spl_,
    g906_n
  );


  or

  (
    g990_n,
    g903_p_spl_,
    g906_p_spl_
  );


  and

  (
    g991_p,
    n2746_lo_p_spl_000,
    lo006_buf_o2_p_spl_00
  );


  or

  (
    g991_n,
    n2746_lo_n_spl_000,
    lo006_buf_o2_n_spl_0
  );


  and

  (
    g992_p,
    g897_n_spl_,
    g900_n_spl_
  );


  or

  (
    g992_n,
    g897_p_spl_,
    g900_p_spl_
  );


  and

  (
    g993_p,
    n2734_lo_p_spl_001,
    lo010_buf_o2_p_spl_00
  );


  or

  (
    g993_n,
    n2734_lo_n_spl_001,
    lo010_buf_o2_n_spl_0
  );


  and

  (
    g994_p,
    n577_o2_p,
    g894_n_spl_
  );


  or

  (
    g994_n,
    n577_o2_n,
    g894_p_spl_
  );


  and

  (
    g995_p,
    n601_o2_n_spl_,
    n625_o2_p_spl_
  );


  or

  (
    g995_n,
    n601_o2_p_spl_,
    n625_o2_n_spl_
  );


  and

  (
    g996_p,
    n601_o2_p_spl_,
    n625_o2_n_spl_
  );


  or

  (
    g996_n,
    n601_o2_n_spl_,
    n625_o2_p_spl_
  );


  and

  (
    g997_p,
    g995_n_spl_,
    g996_n
  );


  or

  (
    g997_n,
    g995_p_spl_,
    g996_p
  );


  and

  (
    g998_p,
    g994_n_spl_,
    g997_p_spl_
  );


  or

  (
    g998_n,
    g994_p_spl_,
    g997_n_spl_
  );


  and

  (
    g999_p,
    g994_p_spl_,
    g997_n_spl_
  );


  or

  (
    g999_n,
    g994_n_spl_,
    g997_p_spl_
  );


  and

  (
    g1000_p,
    g998_n_spl_,
    g999_n
  );


  or

  (
    g1000_n,
    g998_p_spl_,
    g999_p
  );


  and

  (
    g1001_p,
    g993_n_spl_,
    g1000_p_spl_
  );


  or

  (
    g1001_n,
    g993_p_spl_,
    g1000_n_spl_
  );


  and

  (
    g1002_p,
    g993_p_spl_,
    g1000_n_spl_
  );


  or

  (
    g1002_n,
    g993_n_spl_,
    g1000_p_spl_
  );


  and

  (
    g1003_p,
    g1001_n_spl_,
    g1002_n
  );


  or

  (
    g1003_n,
    g1001_p_spl_,
    g1002_p
  );


  and

  (
    g1004_p,
    g992_n_spl_,
    g1003_p_spl_
  );


  or

  (
    g1004_n,
    g992_p_spl_,
    g1003_n_spl_
  );


  and

  (
    g1005_p,
    g992_p_spl_,
    g1003_n_spl_
  );


  or

  (
    g1005_n,
    g992_n_spl_,
    g1003_p_spl_
  );


  and

  (
    g1006_p,
    g1004_n_spl_,
    g1005_n
  );


  or

  (
    g1006_n,
    g1004_p_spl_,
    g1005_p
  );


  and

  (
    g1007_p,
    g991_n_spl_,
    g1006_p_spl_
  );


  or

  (
    g1007_n,
    g991_p_spl_,
    g1006_n_spl_
  );


  and

  (
    g1008_p,
    g991_p_spl_,
    g1006_n_spl_
  );


  or

  (
    g1008_n,
    g991_n_spl_,
    g1006_p_spl_
  );


  and

  (
    g1009_p,
    g1007_n_spl_,
    g1008_n
  );


  or

  (
    g1009_n,
    g1007_p_spl_,
    g1008_p
  );


  and

  (
    g1010_p,
    g990_n_spl_,
    g1009_p_spl_
  );


  or

  (
    g1010_n,
    g990_p_spl_,
    g1009_n_spl_
  );


  and

  (
    g1011_p,
    g990_p_spl_,
    g1009_n_spl_
  );


  or

  (
    g1011_n,
    g990_n_spl_,
    g1009_p_spl_
  );


  and

  (
    g1012_p,
    g1010_n_spl_,
    g1011_n
  );


  or

  (
    g1012_n,
    g1010_p_spl_,
    g1011_p
  );


  or

  (
    g1013_n,
    g887_p,
    g959_p_spl_
  );


  or

  (
    g1014_n,
    g947_n,
    g957_p
  );


  and

  (
    g1015_p,
    g958_n_spl_,
    g1014_n
  );


  and

  (
    g1016_p,
    G1_p_spl_0,
    G19_p_spl_000
  );


  or

  (
    g1016_n,
    G1_n_spl_0,
    G19_n_spl_000
  );


  and

  (
    g1017_p,
    n1808_o2_p,
    n1811_o2_n_spl_
  );


  or

  (
    g1017_n,
    n1808_o2_n,
    n1811_o2_p_spl_
  );


  and

  (
    g1018_p,
    n6036_o2_p_spl_00,
    lo094_buf_o2_p_spl_
  );


  or

  (
    g1018_n,
    n6036_o2_n_spl_0,
    lo094_buf_o2_n_spl_
  );


  and

  (
    g1019_p,
    n1889_o2_p_spl_,
    n1890_o2_n
  );


  or

  (
    g1019_n,
    n1889_o2_n_spl_,
    n1890_o2_p
  );


  and

  (
    g1020_p,
    g1018_n_spl_,
    g1019_p_spl_
  );


  or

  (
    g1020_n,
    g1018_p_spl_,
    g1019_n_spl_
  );


  and

  (
    g1021_p,
    g1018_p_spl_,
    g1019_n_spl_
  );


  or

  (
    g1021_n,
    g1018_n_spl_,
    g1019_p_spl_
  );


  and

  (
    g1022_p,
    g1020_n_spl_,
    g1021_n
  );


  or

  (
    g1022_n,
    g1020_p_spl_,
    g1021_p
  );


  and

  (
    g1023_p,
    g1017_n_spl_,
    g1022_p_spl_
  );


  or

  (
    g1023_n,
    g1017_p_spl_,
    g1022_n_spl_
  );


  and

  (
    g1024_p,
    n6035_o2_p_spl_0,
    lo098_buf_o2_p_spl_00
  );


  or

  (
    g1024_n,
    n6035_o2_n_spl_0,
    lo098_buf_o2_n_spl_00
  );


  and

  (
    g1025_p,
    g1017_p_spl_,
    g1022_n_spl_
  );


  or

  (
    g1025_n,
    g1017_n_spl_,
    g1022_p_spl_
  );


  and

  (
    g1026_p,
    g1023_n_spl_,
    g1025_n
  );


  or

  (
    g1026_n,
    g1023_p_spl_,
    g1025_p
  );


  and

  (
    g1027_p,
    g1024_n_spl_,
    g1026_p_spl_
  );


  or

  (
    g1027_n,
    g1024_p_spl_,
    g1026_n_spl_
  );


  and

  (
    g1028_p,
    g1023_n_spl_,
    g1027_n_spl_
  );


  or

  (
    g1028_n,
    g1023_p_spl_,
    g1027_p_spl_
  );


  and

  (
    g1029_p,
    n6036_o2_p_spl_00,
    lo098_buf_o2_p_spl_00
  );


  or

  (
    g1029_n,
    n6036_o2_n_spl_0,
    lo098_buf_o2_n_spl_00
  );


  and

  (
    g1030_p,
    n6037_o2_p_spl_0,
    lo094_buf_o2_p_spl_
  );


  or

  (
    g1030_n,
    n6037_o2_n_spl_0,
    lo094_buf_o2_n_spl_
  );


  and

  (
    g1031_p,
    n1889_o2_p_spl_,
    g1020_n_spl_
  );


  or

  (
    g1031_n,
    n1889_o2_n_spl_,
    g1020_p_spl_
  );


  and

  (
    g1032_p,
    g1030_n_spl_,
    g1031_n_spl_
  );


  or

  (
    g1032_n,
    g1030_p_spl_,
    g1031_p_spl_
  );


  and

  (
    g1033_p,
    g1030_p_spl_,
    g1031_p_spl_
  );


  or

  (
    g1033_n,
    g1030_n_spl_,
    g1031_n_spl_
  );


  and

  (
    g1034_p,
    g1032_n_spl_,
    g1033_n
  );


  or

  (
    g1034_n,
    g1032_p_spl_,
    g1033_p
  );


  and

  (
    g1035_p,
    g1029_n_spl_,
    g1034_p_spl_
  );


  or

  (
    g1035_n,
    g1029_p_spl_,
    g1034_n_spl_
  );


  and

  (
    g1036_p,
    g1029_p_spl_,
    g1034_n_spl_
  );


  or

  (
    g1036_n,
    g1029_n_spl_,
    g1034_p_spl_
  );


  and

  (
    g1037_p,
    g1035_n_spl_,
    g1036_n
  );


  or

  (
    g1037_n,
    g1035_p_spl_,
    g1036_p
  );


  and

  (
    g1038_p,
    g1028_n_spl_,
    g1037_p_spl_
  );


  or

  (
    g1038_n,
    g1028_p_spl_,
    g1037_n_spl_
  );


  and

  (
    g1039_p,
    n6035_o2_p_spl_0,
    lo102_buf_o2_p_spl_010
  );


  or

  (
    g1039_n,
    n6035_o2_n_spl_0,
    lo102_buf_o2_n_spl_010
  );


  and

  (
    g1040_p,
    g1028_p_spl_,
    g1037_n_spl_
  );


  or

  (
    g1040_n,
    g1028_n_spl_,
    g1037_p_spl_
  );


  and

  (
    g1041_p,
    g1038_n_spl_,
    g1040_n
  );


  or

  (
    g1041_n,
    g1038_p_spl_,
    g1040_p
  );


  and

  (
    g1042_p,
    g1039_n_spl_,
    g1041_p_spl_
  );


  or

  (
    g1042_n,
    g1039_p_spl_,
    g1041_n_spl_
  );


  and

  (
    g1043_p,
    g1038_n_spl_,
    g1042_n_spl_
  );


  or

  (
    g1043_n,
    g1038_p_spl_,
    g1042_p_spl_
  );


  and

  (
    g1044_p,
    n6036_o2_p_spl_0,
    lo102_buf_o2_p_spl_010
  );


  or

  (
    g1044_n,
    n6036_o2_n_spl_,
    lo102_buf_o2_n_spl_010
  );


  and

  (
    g1045_p,
    n6037_o2_p_spl_0,
    lo098_buf_o2_p_spl_0
  );


  or

  (
    g1045_n,
    n6037_o2_n_spl_0,
    lo098_buf_o2_n_spl_0
  );


  and

  (
    g1046_p,
    g1032_n_spl_,
    g1035_n_spl_
  );


  or

  (
    g1046_n,
    g1032_p_spl_,
    g1035_p_spl_
  );


  and

  (
    g1047_p,
    g1045_n_spl_,
    g1046_n_spl_
  );


  or

  (
    g1047_n,
    g1045_p_spl_,
    g1046_p_spl_
  );


  and

  (
    g1048_p,
    g1045_p_spl_,
    g1046_p_spl_
  );


  or

  (
    g1048_n,
    g1045_n_spl_,
    g1046_n_spl_
  );


  and

  (
    g1049_p,
    g1047_n_spl_,
    g1048_n
  );


  or

  (
    g1049_n,
    g1047_p_spl_,
    g1048_p
  );


  and

  (
    g1050_p,
    g1044_n_spl_,
    g1049_p_spl_
  );


  or

  (
    g1050_n,
    g1044_p_spl_,
    g1049_n_spl_
  );


  and

  (
    g1051_p,
    g1044_p_spl_,
    g1049_n_spl_
  );


  or

  (
    g1051_n,
    g1044_n_spl_,
    g1049_p_spl_
  );


  and

  (
    g1052_p,
    g1050_n_spl_,
    g1051_n
  );


  or

  (
    g1052_n,
    g1050_p_spl_,
    g1051_p
  );


  and

  (
    g1053_p,
    g1043_n_spl_,
    g1052_p_spl_
  );


  or

  (
    g1053_n,
    g1043_p_spl_,
    g1052_n_spl_
  );


  and

  (
    g1054_p,
    n1628_o2_p,
    n1631_o2_n_spl_
  );


  or

  (
    g1054_n,
    n1628_o2_n,
    n1631_o2_p_spl_
  );


  and

  (
    g1055_p,
    n6033_o2_p_spl_00,
    lo098_buf_o2_p_spl_1
  );


  or

  (
    g1055_n,
    n6033_o2_n_spl_0,
    lo098_buf_o2_n_spl_1
  );


  and

  (
    g1056_p,
    n1725_o2_p_spl_,
    n1726_o2_n
  );


  or

  (
    g1056_n,
    n1725_o2_n_spl_,
    n1726_o2_p
  );


  and

  (
    g1057_p,
    g1055_n_spl_,
    g1056_p_spl_
  );


  or

  (
    g1057_n,
    g1055_p_spl_,
    g1056_n_spl_
  );


  and

  (
    g1058_p,
    g1055_p_spl_,
    g1056_n_spl_
  );


  or

  (
    g1058_n,
    g1055_n_spl_,
    g1056_p_spl_
  );


  and

  (
    g1059_p,
    g1057_n_spl_,
    g1058_n
  );


  or

  (
    g1059_n,
    g1057_p_spl_,
    g1058_p
  );


  and

  (
    g1060_p,
    g1054_n_spl_,
    g1059_p_spl_
  );


  or

  (
    g1060_n,
    g1054_p_spl_,
    g1059_n_spl_
  );


  and

  (
    g1061_p,
    n6032_o2_p_spl_0,
    lo102_buf_o2_p_spl_011
  );


  or

  (
    g1061_n,
    n6032_o2_n_spl_0,
    lo102_buf_o2_n_spl_011
  );


  and

  (
    g1062_p,
    g1054_p_spl_,
    g1059_n_spl_
  );


  or

  (
    g1062_n,
    g1054_n_spl_,
    g1059_p_spl_
  );


  and

  (
    g1063_p,
    g1060_n_spl_,
    g1062_n
  );


  or

  (
    g1063_n,
    g1060_p_spl_,
    g1062_p
  );


  and

  (
    g1064_p,
    g1061_n_spl_,
    g1063_p_spl_
  );


  or

  (
    g1064_n,
    g1061_p_spl_,
    g1063_n_spl_
  );


  and

  (
    g1065_p,
    g1060_n_spl_,
    g1064_n_spl_
  );


  or

  (
    g1065_n,
    g1060_p_spl_,
    g1064_p_spl_
  );


  and

  (
    g1066_p,
    n6033_o2_p_spl_00,
    lo102_buf_o2_p_spl_011
  );


  or

  (
    g1066_n,
    n6033_o2_n_spl_0,
    lo102_buf_o2_n_spl_011
  );


  and

  (
    g1067_p,
    n1725_o2_p_spl_,
    g1057_n_spl_
  );


  or

  (
    g1067_n,
    n1725_o2_n_spl_,
    g1057_p_spl_
  );


  and

  (
    g1068_p,
    n6034_o2_p_spl_0,
    lo098_buf_o2_p_spl_1
  );


  or

  (
    g1068_n,
    n6034_o2_n_spl_0,
    lo098_buf_o2_n_spl_1
  );


  and

  (
    g1069_p,
    n1719_o2_p,
    n1722_o2_n
  );


  or

  (
    g1069_n,
    n1719_o2_n,
    n1722_o2_p
  );


  and

  (
    g1070_p,
    n1811_o2_n_spl_,
    n1812_o2_n
  );


  or

  (
    g1070_n,
    n1811_o2_p_spl_,
    n1812_o2_p
  );


  and

  (
    g1071_p,
    g1069_n_spl_,
    g1070_p_spl_
  );


  or

  (
    g1071_n,
    g1069_p_spl_,
    g1070_n_spl_
  );


  and

  (
    g1072_p,
    g1069_p_spl_,
    g1070_n_spl_
  );


  or

  (
    g1072_n,
    g1069_n_spl_,
    g1070_p_spl_
  );


  and

  (
    g1073_p,
    g1071_n_spl_,
    g1072_n
  );


  or

  (
    g1073_n,
    g1071_p_spl_,
    g1072_p
  );


  and

  (
    g1074_p,
    g1068_n_spl_,
    g1073_p_spl_
  );


  or

  (
    g1074_n,
    g1068_p_spl_,
    g1073_n_spl_
  );


  and

  (
    g1075_p,
    g1068_p_spl_,
    g1073_n_spl_
  );


  or

  (
    g1075_n,
    g1068_n_spl_,
    g1073_p_spl_
  );


  and

  (
    g1076_p,
    g1074_n_spl_,
    g1075_n
  );


  or

  (
    g1076_n,
    g1074_p_spl_,
    g1075_p
  );


  and

  (
    g1077_p,
    g1067_n_spl_,
    g1076_p_spl_
  );


  or

  (
    g1077_n,
    g1067_p_spl_,
    g1076_n_spl_
  );


  and

  (
    g1078_p,
    g1067_p_spl_,
    g1076_n_spl_
  );


  or

  (
    g1078_n,
    g1067_n_spl_,
    g1076_p_spl_
  );


  and

  (
    g1079_p,
    g1077_n_spl_,
    g1078_n
  );


  or

  (
    g1079_n,
    g1077_p_spl_,
    g1078_p
  );


  and

  (
    g1080_p,
    g1066_n_spl_,
    g1079_p_spl_
  );


  or

  (
    g1080_n,
    g1066_p_spl_,
    g1079_n_spl_
  );


  and

  (
    g1081_p,
    g1066_p_spl_,
    g1079_n_spl_
  );


  or

  (
    g1081_n,
    g1066_n_spl_,
    g1079_p_spl_
  );


  and

  (
    g1082_p,
    g1080_n_spl_,
    g1081_n
  );


  or

  (
    g1082_n,
    g1080_p_spl_,
    g1081_p
  );


  and

  (
    g1083_p,
    g1065_n_spl_,
    g1082_p_spl_
  );


  or

  (
    g1083_n,
    g1065_p_spl_,
    g1082_n_spl_
  );


  and

  (
    g1084_p,
    n2797_lo_p_spl_001,
    n6032_o2_p_spl_0
  );


  or

  (
    g1084_n,
    n2797_lo_n_spl_001,
    n6032_o2_n_spl_0
  );


  and

  (
    g1085_p,
    g1065_p_spl_,
    g1082_n_spl_
  );


  or

  (
    g1085_n,
    g1065_n_spl_,
    g1082_p_spl_
  );


  and

  (
    g1086_p,
    g1083_n_spl_,
    g1085_n
  );


  or

  (
    g1086_n,
    g1083_p_spl_,
    g1085_p
  );


  and

  (
    g1087_p,
    g1084_n_spl_,
    g1086_p_spl_
  );


  or

  (
    g1087_n,
    g1084_p_spl_,
    g1086_n_spl_
  );


  and

  (
    g1088_p,
    g1083_n_spl_,
    g1087_n_spl_
  );


  or

  (
    g1088_n,
    g1083_p_spl_,
    g1087_p_spl_
  );


  and

  (
    g1089_p,
    n2797_lo_p_spl_010,
    n6033_o2_p_spl_0
  );


  or

  (
    g1089_n,
    n2797_lo_n_spl_010,
    n6033_o2_n_spl_
  );


  and

  (
    g1090_p,
    g1077_n_spl_,
    g1080_n_spl_
  );


  or

  (
    g1090_n,
    g1077_p_spl_,
    g1080_p_spl_
  );


  and

  (
    g1091_p,
    n6034_o2_p_spl_0,
    lo102_buf_o2_p_spl_100
  );


  or

  (
    g1091_n,
    n6034_o2_n_spl_0,
    lo102_buf_o2_n_spl_100
  );


  and

  (
    g1092_p,
    g1071_n_spl_,
    g1074_n_spl_
  );


  or

  (
    g1092_n,
    g1071_p_spl_,
    g1074_p_spl_
  );


  and

  (
    g1093_p,
    g1024_p_spl_,
    g1026_n_spl_
  );


  or

  (
    g1093_n,
    g1024_n_spl_,
    g1026_p_spl_
  );


  and

  (
    g1094_p,
    g1027_n_spl_,
    g1093_n
  );


  or

  (
    g1094_n,
    g1027_p_spl_,
    g1093_p
  );


  and

  (
    g1095_p,
    g1092_n_spl_,
    g1094_p_spl_
  );


  or

  (
    g1095_n,
    g1092_p_spl_,
    g1094_n_spl_
  );


  and

  (
    g1096_p,
    g1092_p_spl_,
    g1094_n_spl_
  );


  or

  (
    g1096_n,
    g1092_n_spl_,
    g1094_p_spl_
  );


  and

  (
    g1097_p,
    g1095_n_spl_,
    g1096_n
  );


  or

  (
    g1097_n,
    g1095_p_spl_,
    g1096_p
  );


  and

  (
    g1098_p,
    g1091_n_spl_,
    g1097_p_spl_
  );


  or

  (
    g1098_n,
    g1091_p_spl_,
    g1097_n_spl_
  );


  and

  (
    g1099_p,
    g1091_p_spl_,
    g1097_n_spl_
  );


  or

  (
    g1099_n,
    g1091_n_spl_,
    g1097_p_spl_
  );


  and

  (
    g1100_p,
    g1098_n_spl_,
    g1099_n
  );


  or

  (
    g1100_n,
    g1098_p_spl_,
    g1099_p
  );


  and

  (
    g1101_p,
    g1090_n_spl_,
    g1100_p_spl_
  );


  or

  (
    g1101_n,
    g1090_p_spl_,
    g1100_n_spl_
  );


  and

  (
    g1102_p,
    g1090_p_spl_,
    g1100_n_spl_
  );


  or

  (
    g1102_n,
    g1090_n_spl_,
    g1100_p_spl_
  );


  and

  (
    g1103_p,
    g1101_n_spl_,
    g1102_n
  );


  or

  (
    g1103_n,
    g1101_p_spl_,
    g1102_p
  );


  and

  (
    g1104_p,
    g1089_n_spl_,
    g1103_p_spl_
  );


  or

  (
    g1104_n,
    g1089_p_spl_,
    g1103_n_spl_
  );


  and

  (
    g1105_p,
    g1089_p_spl_,
    g1103_n_spl_
  );


  or

  (
    g1105_n,
    g1089_n_spl_,
    g1103_p_spl_
  );


  and

  (
    g1106_p,
    g1104_n_spl_,
    g1105_n
  );


  or

  (
    g1106_n,
    g1104_p_spl_,
    g1105_p
  );


  and

  (
    g1107_p,
    g1088_n_spl_,
    g1106_p_spl_
  );


  or

  (
    g1107_n,
    g1088_p_spl_,
    g1106_n_spl_
  );


  and

  (
    g1108_p,
    n6029_o2_p_spl_00,
    lo102_buf_o2_p_spl_100
  );


  or

  (
    g1108_n,
    n6029_o2_n_spl_0,
    lo102_buf_o2_n_spl_100
  );


  and

  (
    g1109_p,
    n1420_o2_p_spl_,
    n1421_o2_n
  );


  or

  (
    g1109_n,
    n1420_o2_n_spl_,
    n1421_o2_p
  );


  and

  (
    g1110_p,
    g1108_n_spl_,
    g1109_p_spl_
  );


  or

  (
    g1110_n,
    g1108_p_spl_,
    g1109_n_spl_
  );


  and

  (
    g1111_p,
    n1420_o2_p_spl_,
    g1110_n_spl_
  );


  or

  (
    g1111_n,
    n1420_o2_n_spl_,
    g1110_p_spl_
  );


  and

  (
    g1112_p,
    n6030_o2_p_spl_00,
    lo102_buf_o2_p_spl_101
  );


  or

  (
    g1112_n,
    n6030_o2_n_spl_0,
    lo102_buf_o2_n_spl_101
  );


  and

  (
    g1113_p,
    n1529_o2_p_spl_,
    n1530_o2_n
  );


  or

  (
    g1113_n,
    n1529_o2_n_spl_,
    n1530_o2_p
  );


  and

  (
    g1114_p,
    g1112_n_spl_,
    g1113_p_spl_
  );


  or

  (
    g1114_n,
    g1112_p_spl_,
    g1113_n_spl_
  );


  and

  (
    g1115_p,
    g1112_p_spl_,
    g1113_n_spl_
  );


  or

  (
    g1115_n,
    g1112_n_spl_,
    g1113_p_spl_
  );


  and

  (
    g1116_p,
    g1114_n_spl_,
    g1115_n
  );


  or

  (
    g1116_n,
    g1114_p_spl_,
    g1115_p
  );


  and

  (
    g1117_p,
    g1111_n_spl_,
    g1116_p_spl_
  );


  or

  (
    g1117_n,
    g1111_p_spl_,
    g1116_n_spl_
  );


  and

  (
    g1118_p,
    n2797_lo_p_spl_010,
    n6029_o2_p_spl_00
  );


  or

  (
    g1118_n,
    n2797_lo_n_spl_010,
    n6029_o2_n_spl_0
  );


  and

  (
    g1119_p,
    g1111_p_spl_,
    g1116_n_spl_
  );


  or

  (
    g1119_n,
    g1111_n_spl_,
    g1116_p_spl_
  );


  and

  (
    g1120_p,
    g1117_n_spl_,
    g1119_n
  );


  or

  (
    g1120_n,
    g1117_p_spl_,
    g1119_p
  );


  and

  (
    g1121_p,
    g1118_n_spl_,
    g1120_p_spl_
  );


  or

  (
    g1121_n,
    g1118_p_spl_,
    g1120_n_spl_
  );


  and

  (
    g1122_p,
    g1117_n_spl_,
    g1121_n_spl_
  );


  or

  (
    g1122_n,
    g1117_p_spl_,
    g1121_p_spl_
  );


  and

  (
    g1123_p,
    n2797_lo_p_spl_011,
    n6030_o2_p_spl_00
  );


  or

  (
    g1123_n,
    n2797_lo_n_spl_011,
    n6030_o2_n_spl_0
  );


  and

  (
    g1124_p,
    n1529_o2_p_spl_,
    g1114_n_spl_
  );


  or

  (
    g1124_n,
    n1529_o2_n_spl_,
    g1114_p_spl_
  );


  and

  (
    g1125_p,
    n6031_o2_p_spl_0,
    lo102_buf_o2_p_spl_101
  );


  or

  (
    g1125_n,
    n6031_o2_n_spl_0,
    lo102_buf_o2_n_spl_101
  );


  and

  (
    g1126_p,
    n1523_o2_p,
    n1526_o2_n
  );


  or

  (
    g1126_n,
    n1523_o2_n,
    n1526_o2_p
  );


  and

  (
    g1127_p,
    n1631_o2_n_spl_,
    n1632_o2_n
  );


  or

  (
    g1127_n,
    n1631_o2_p_spl_,
    n1632_o2_p
  );


  and

  (
    g1128_p,
    g1126_n_spl_,
    g1127_p_spl_
  );


  or

  (
    g1128_n,
    g1126_p_spl_,
    g1127_n_spl_
  );


  and

  (
    g1129_p,
    g1126_p_spl_,
    g1127_n_spl_
  );


  or

  (
    g1129_n,
    g1126_n_spl_,
    g1127_p_spl_
  );


  and

  (
    g1130_p,
    g1128_n_spl_,
    g1129_n
  );


  or

  (
    g1130_n,
    g1128_p_spl_,
    g1129_p
  );


  and

  (
    g1131_p,
    g1125_n_spl_,
    g1130_p_spl_
  );


  or

  (
    g1131_n,
    g1125_p_spl_,
    g1130_n_spl_
  );


  and

  (
    g1132_p,
    g1125_p_spl_,
    g1130_n_spl_
  );


  or

  (
    g1132_n,
    g1125_n_spl_,
    g1130_p_spl_
  );


  and

  (
    g1133_p,
    g1131_n_spl_,
    g1132_n
  );


  or

  (
    g1133_n,
    g1131_p_spl_,
    g1132_p
  );


  and

  (
    g1134_p,
    g1124_n_spl_,
    g1133_p_spl_
  );


  or

  (
    g1134_n,
    g1124_p_spl_,
    g1133_n_spl_
  );


  and

  (
    g1135_p,
    g1124_p_spl_,
    g1133_n_spl_
  );


  or

  (
    g1135_n,
    g1124_n_spl_,
    g1133_p_spl_
  );


  and

  (
    g1136_p,
    g1134_n_spl_,
    g1135_n
  );


  or

  (
    g1136_n,
    g1134_p_spl_,
    g1135_p
  );


  and

  (
    g1137_p,
    g1123_n_spl_,
    g1136_p_spl_
  );


  or

  (
    g1137_n,
    g1123_p_spl_,
    g1136_n_spl_
  );


  and

  (
    g1138_p,
    g1123_p_spl_,
    g1136_n_spl_
  );


  or

  (
    g1138_n,
    g1123_n_spl_,
    g1136_p_spl_
  );


  and

  (
    g1139_p,
    g1137_n_spl_,
    g1138_n
  );


  or

  (
    g1139_n,
    g1137_p_spl_,
    g1138_p
  );


  and

  (
    g1140_p,
    g1122_n_spl_,
    g1139_p_spl_
  );


  or

  (
    g1140_n,
    g1122_p_spl_,
    g1139_n_spl_
  );


  and

  (
    g1141_p,
    n2809_lo_p_spl_001,
    n6029_o2_p_spl_0
  );


  or

  (
    g1141_n,
    n2809_lo_n_spl_001,
    n6029_o2_n_spl_1
  );


  and

  (
    g1142_p,
    g1122_p_spl_,
    g1139_n_spl_
  );


  or

  (
    g1142_n,
    g1122_n_spl_,
    g1139_p_spl_
  );


  and

  (
    g1143_p,
    g1140_n_spl_,
    g1142_n
  );


  or

  (
    g1143_n,
    g1140_p_spl_,
    g1142_p
  );


  and

  (
    g1144_p,
    g1141_n_spl_,
    g1143_p_spl_
  );


  or

  (
    g1144_n,
    g1141_p_spl_,
    g1143_n_spl_
  );


  and

  (
    g1145_p,
    g1140_n_spl_,
    g1144_n_spl_
  );


  or

  (
    g1145_n,
    g1140_p_spl_,
    g1144_p_spl_
  );


  and

  (
    g1146_p,
    n2809_lo_p_spl_001,
    n6030_o2_p_spl_0
  );


  or

  (
    g1146_n,
    n2809_lo_n_spl_001,
    n6030_o2_n_spl_
  );


  and

  (
    g1147_p,
    g1134_n_spl_,
    g1137_n_spl_
  );


  or

  (
    g1147_n,
    g1134_p_spl_,
    g1137_p_spl_
  );


  and

  (
    g1148_p,
    n2797_lo_p_spl_011,
    n6031_o2_p_spl_0
  );


  or

  (
    g1148_n,
    n2797_lo_n_spl_011,
    n6031_o2_n_spl_0
  );


  and

  (
    g1149_p,
    g1128_n_spl_,
    g1131_n_spl_
  );


  or

  (
    g1149_n,
    g1128_p_spl_,
    g1131_p_spl_
  );


  and

  (
    g1150_p,
    g1061_p_spl_,
    g1063_n_spl_
  );


  or

  (
    g1150_n,
    g1061_n_spl_,
    g1063_p_spl_
  );


  and

  (
    g1151_p,
    g1064_n_spl_,
    g1150_n
  );


  or

  (
    g1151_n,
    g1064_p_spl_,
    g1150_p
  );


  and

  (
    g1152_p,
    g1149_n_spl_,
    g1151_p_spl_
  );


  or

  (
    g1152_n,
    g1149_p_spl_,
    g1151_n_spl_
  );


  and

  (
    g1153_p,
    g1149_p_spl_,
    g1151_n_spl_
  );


  or

  (
    g1153_n,
    g1149_n_spl_,
    g1151_p_spl_
  );


  and

  (
    g1154_p,
    g1152_n_spl_,
    g1153_n
  );


  or

  (
    g1154_n,
    g1152_p_spl_,
    g1153_p
  );


  and

  (
    g1155_p,
    g1148_n_spl_,
    g1154_p_spl_
  );


  or

  (
    g1155_n,
    g1148_p_spl_,
    g1154_n_spl_
  );


  and

  (
    g1156_p,
    g1148_p_spl_,
    g1154_n_spl_
  );


  or

  (
    g1156_n,
    g1148_n_spl_,
    g1154_p_spl_
  );


  and

  (
    g1157_p,
    g1155_n_spl_,
    g1156_n
  );


  or

  (
    g1157_n,
    g1155_p_spl_,
    g1156_p
  );


  and

  (
    g1158_p,
    g1147_n_spl_,
    g1157_p_spl_
  );


  or

  (
    g1158_n,
    g1147_p_spl_,
    g1157_n_spl_
  );


  and

  (
    g1159_p,
    g1147_p_spl_,
    g1157_n_spl_
  );


  or

  (
    g1159_n,
    g1147_n_spl_,
    g1157_p_spl_
  );


  and

  (
    g1160_p,
    g1158_n_spl_,
    g1159_n
  );


  or

  (
    g1160_n,
    g1158_p_spl_,
    g1159_p
  );


  and

  (
    g1161_p,
    g1146_n_spl_,
    g1160_p_spl_
  );


  or

  (
    g1161_n,
    g1146_p_spl_,
    g1160_n_spl_
  );


  and

  (
    g1162_p,
    g1146_p_spl_,
    g1160_n_spl_
  );


  or

  (
    g1162_n,
    g1146_n_spl_,
    g1160_p_spl_
  );


  and

  (
    g1163_p,
    g1161_n_spl_,
    g1162_n
  );


  or

  (
    g1163_n,
    g1161_p_spl_,
    g1162_p
  );


  and

  (
    g1164_p,
    g1145_n_spl_,
    g1163_p_spl_
  );


  or

  (
    g1164_n,
    g1145_p_spl_,
    g1163_n_spl_
  );


  and

  (
    g1165_p,
    n6026_o2_p_spl_00,
    lo102_buf_o2_p_spl_110
  );


  or

  (
    g1165_n,
    n6026_o2_n_spl_00,
    lo102_buf_o2_n_spl_110
  );


  and

  (
    g1166_p,
    n1097_o2_p_spl_,
    n1098_o2_n
  );


  or

  (
    g1166_n,
    n1097_o2_n_spl_,
    n1098_o2_p
  );


  and

  (
    g1167_p,
    g1165_n_spl_,
    g1166_p_spl_
  );


  or

  (
    g1167_n,
    g1165_p_spl_,
    g1166_n_spl_
  );


  and

  (
    g1168_p,
    n1097_o2_p_spl_,
    g1167_n_spl_
  );


  or

  (
    g1168_n,
    n1097_o2_n_spl_,
    g1167_p_spl_
  );


  and

  (
    g1169_p,
    n6027_o2_p_spl_00,
    lo102_buf_o2_p_spl_110
  );


  or

  (
    g1169_n,
    n6027_o2_n_spl_0,
    lo102_buf_o2_n_spl_110
  );


  and

  (
    g1170_p,
    n1199_o2_p_spl_,
    n1200_o2_n
  );


  or

  (
    g1170_n,
    n1199_o2_n_spl_,
    n1200_o2_p
  );


  and

  (
    g1171_p,
    g1169_n_spl_,
    g1170_p_spl_
  );


  or

  (
    g1171_n,
    g1169_p_spl_,
    g1170_n_spl_
  );


  and

  (
    g1172_p,
    g1169_p_spl_,
    g1170_n_spl_
  );


  or

  (
    g1172_n,
    g1169_n_spl_,
    g1170_p_spl_
  );


  and

  (
    g1173_p,
    g1171_n_spl_,
    g1172_n
  );


  or

  (
    g1173_n,
    g1171_p_spl_,
    g1172_p
  );


  and

  (
    g1174_p,
    g1168_n_spl_,
    g1173_p_spl_
  );


  or

  (
    g1174_n,
    g1168_p_spl_,
    g1173_n_spl_
  );


  and

  (
    g1175_p,
    n2797_lo_p_spl_100,
    n6026_o2_p_spl_00
  );


  or

  (
    g1175_n,
    n2797_lo_n_spl_100,
    n6026_o2_n_spl_00
  );


  and

  (
    g1176_p,
    g1168_p_spl_,
    g1173_n_spl_
  );


  or

  (
    g1176_n,
    g1168_n_spl_,
    g1173_p_spl_
  );


  and

  (
    g1177_p,
    g1174_n_spl_,
    g1176_n
  );


  or

  (
    g1177_n,
    g1174_p_spl_,
    g1176_p
  );


  and

  (
    g1178_p,
    g1175_n_spl_,
    g1177_p_spl_
  );


  or

  (
    g1178_n,
    g1175_p_spl_,
    g1177_n_spl_
  );


  and

  (
    g1179_p,
    g1174_n_spl_,
    g1178_n_spl_
  );


  or

  (
    g1179_n,
    g1174_p_spl_,
    g1178_p_spl_
  );


  and

  (
    g1180_p,
    n2797_lo_p_spl_100,
    n6027_o2_p_spl_00
  );


  or

  (
    g1180_n,
    n2797_lo_n_spl_100,
    n6027_o2_n_spl_0
  );


  and

  (
    g1181_p,
    n1199_o2_p_spl_,
    g1171_n_spl_
  );


  or

  (
    g1181_n,
    n1199_o2_n_spl_,
    g1171_p_spl_
  );


  and

  (
    g1182_p,
    n6028_o2_p_spl_00,
    lo102_buf_o2_p_spl_111
  );


  or

  (
    g1182_n,
    n6028_o2_n_spl_0,
    lo102_buf_o2_n_spl_111
  );


  and

  (
    g1183_p,
    n1309_o2_p_spl_,
    n1310_o2_n
  );


  or

  (
    g1183_n,
    n1309_o2_n_spl_,
    n1310_o2_p
  );


  and

  (
    g1184_p,
    g1182_n_spl_,
    g1183_p_spl_
  );


  or

  (
    g1184_n,
    g1182_p_spl_,
    g1183_n_spl_
  );


  and

  (
    g1185_p,
    g1182_p_spl_,
    g1183_n_spl_
  );


  or

  (
    g1185_n,
    g1182_n_spl_,
    g1183_p_spl_
  );


  and

  (
    g1186_p,
    g1184_n_spl_,
    g1185_n
  );


  or

  (
    g1186_n,
    g1184_p_spl_,
    g1185_p
  );


  and

  (
    g1187_p,
    g1181_n_spl_,
    g1186_p_spl_
  );


  or

  (
    g1187_n,
    g1181_p_spl_,
    g1186_n_spl_
  );


  and

  (
    g1188_p,
    g1181_p_spl_,
    g1186_n_spl_
  );


  or

  (
    g1188_n,
    g1181_n_spl_,
    g1186_p_spl_
  );


  and

  (
    g1189_p,
    g1187_n_spl_,
    g1188_n
  );


  or

  (
    g1189_n,
    g1187_p_spl_,
    g1188_p
  );


  and

  (
    g1190_p,
    g1180_n_spl_,
    g1189_p_spl_
  );


  or

  (
    g1190_n,
    g1180_p_spl_,
    g1189_n_spl_
  );


  and

  (
    g1191_p,
    g1180_p_spl_,
    g1189_n_spl_
  );


  or

  (
    g1191_n,
    g1180_n_spl_,
    g1189_p_spl_
  );


  and

  (
    g1192_p,
    g1190_n_spl_,
    g1191_n
  );


  or

  (
    g1192_n,
    g1190_p_spl_,
    g1191_p
  );


  and

  (
    g1193_p,
    g1179_n_spl_,
    g1192_p_spl_
  );


  or

  (
    g1193_n,
    g1179_p_spl_,
    g1192_n_spl_
  );


  and

  (
    g1194_p,
    n2809_lo_p_spl_010,
    n6026_o2_p_spl_01
  );


  or

  (
    g1194_n,
    n2809_lo_n_spl_010,
    n6026_o2_n_spl_0
  );


  and

  (
    g1195_p,
    g1179_p_spl_,
    g1192_n_spl_
  );


  or

  (
    g1195_n,
    g1179_n_spl_,
    g1192_p_spl_
  );


  and

  (
    g1196_p,
    g1193_n_spl_,
    g1195_n
  );


  or

  (
    g1196_n,
    g1193_p_spl_,
    g1195_p
  );


  and

  (
    g1197_p,
    g1194_n_spl_,
    g1196_p_spl_
  );


  or

  (
    g1197_n,
    g1194_p_spl_,
    g1196_n_spl_
  );


  and

  (
    g1198_p,
    g1193_n_spl_,
    g1197_n_spl_
  );


  or

  (
    g1198_n,
    g1193_p_spl_,
    g1197_p_spl_
  );


  and

  (
    g1199_p,
    n2809_lo_p_spl_010,
    n6027_o2_p_spl_01
  );


  or

  (
    g1199_n,
    n2809_lo_n_spl_010,
    n6027_o2_n_spl_1
  );


  and

  (
    g1200_p,
    g1187_n_spl_,
    g1190_n_spl_
  );


  or

  (
    g1200_n,
    g1187_p_spl_,
    g1190_p_spl_
  );


  and

  (
    g1201_p,
    n2797_lo_p_spl_101,
    n6028_o2_p_spl_00
  );


  or

  (
    g1201_n,
    n2797_lo_n_spl_101,
    n6028_o2_n_spl_0
  );


  and

  (
    g1202_p,
    n1309_o2_p_spl_,
    g1184_n_spl_
  );


  or

  (
    g1202_n,
    n1309_o2_n_spl_,
    g1184_p_spl_
  );


  and

  (
    g1203_p,
    g1108_p_spl_,
    g1109_n_spl_
  );


  or

  (
    g1203_n,
    g1108_n_spl_,
    g1109_p_spl_
  );


  and

  (
    g1204_p,
    g1110_n_spl_,
    g1203_n
  );


  or

  (
    g1204_n,
    g1110_p_spl_,
    g1203_p
  );


  and

  (
    g1205_p,
    g1202_n_spl_,
    g1204_p_spl_
  );


  or

  (
    g1205_n,
    g1202_p_spl_,
    g1204_n_spl_
  );


  and

  (
    g1206_p,
    g1202_p_spl_,
    g1204_n_spl_
  );


  or

  (
    g1206_n,
    g1202_n_spl_,
    g1204_p_spl_
  );


  and

  (
    g1207_p,
    g1205_n_spl_,
    g1206_n
  );


  or

  (
    g1207_n,
    g1205_p_spl_,
    g1206_p
  );


  and

  (
    g1208_p,
    g1201_n_spl_,
    g1207_p_spl_
  );


  or

  (
    g1208_n,
    g1201_p_spl_,
    g1207_n_spl_
  );


  and

  (
    g1209_p,
    g1201_p_spl_,
    g1207_n_spl_
  );


  or

  (
    g1209_n,
    g1201_n_spl_,
    g1207_p_spl_
  );


  and

  (
    g1210_p,
    g1208_n_spl_,
    g1209_n
  );


  or

  (
    g1210_n,
    g1208_p_spl_,
    g1209_p
  );


  and

  (
    g1211_p,
    g1200_n_spl_,
    g1210_p_spl_
  );


  or

  (
    g1211_n,
    g1200_p_spl_,
    g1210_n_spl_
  );


  and

  (
    g1212_p,
    g1200_p_spl_,
    g1210_n_spl_
  );


  or

  (
    g1212_n,
    g1200_n_spl_,
    g1210_p_spl_
  );


  and

  (
    g1213_p,
    g1211_n_spl_,
    g1212_n
  );


  or

  (
    g1213_n,
    g1211_p_spl_,
    g1212_p
  );


  and

  (
    g1214_p,
    g1199_n_spl_,
    g1213_p_spl_
  );


  or

  (
    g1214_n,
    g1199_p_spl_,
    g1213_n_spl_
  );


  and

  (
    g1215_p,
    g1199_p_spl_,
    g1213_n_spl_
  );


  or

  (
    g1215_n,
    g1199_n_spl_,
    g1213_p_spl_
  );


  and

  (
    g1216_p,
    g1214_n_spl_,
    g1215_n
  );


  or

  (
    g1216_n,
    g1214_p_spl_,
    g1215_p
  );


  and

  (
    g1217_p,
    g1198_n_spl_,
    g1216_p_spl_
  );


  or

  (
    g1217_n,
    g1198_p_spl_,
    g1216_n_spl_
  );


  and

  (
    g1218_p,
    n2821_lo_p_spl_000,
    n6026_o2_p_spl_01
  );


  or

  (
    g1218_n,
    n2821_lo_n_spl_00,
    n6026_o2_n_spl_1
  );


  and

  (
    g1219_p,
    g1198_p_spl_,
    g1216_n_spl_
  );


  or

  (
    g1219_n,
    g1198_n_spl_,
    g1216_p_spl_
  );


  and

  (
    g1220_p,
    g1217_n_spl_,
    g1219_n
  );


  or

  (
    g1220_n,
    g1217_p_spl_,
    g1219_p
  );


  and

  (
    g1221_p,
    g1218_n_spl_,
    g1220_p_spl_
  );


  or

  (
    g1221_n,
    g1218_p_spl_,
    g1220_n_spl_
  );


  and

  (
    g1222_p,
    g1217_n_spl_,
    g1221_n_spl_
  );


  or

  (
    g1222_n,
    g1217_p_spl_,
    g1221_p_spl_
  );


  and

  (
    g1223_p,
    n2821_lo_p_spl_001,
    n6027_o2_p_spl_01
  );


  or

  (
    g1223_n,
    n2821_lo_n_spl_01,
    n6027_o2_n_spl_1
  );


  and

  (
    g1224_p,
    g1211_n_spl_,
    g1214_n_spl_
  );


  or

  (
    g1224_n,
    g1211_p_spl_,
    g1214_p_spl_
  );


  and

  (
    g1225_p,
    n2809_lo_p_spl_011,
    n6028_o2_p_spl_0
  );


  or

  (
    g1225_n,
    n2809_lo_n_spl_01,
    n6028_o2_n_spl_1
  );


  and

  (
    g1226_p,
    g1205_n_spl_,
    g1208_n_spl_
  );


  or

  (
    g1226_n,
    g1205_p_spl_,
    g1208_p_spl_
  );


  and

  (
    g1227_p,
    g1118_p_spl_,
    g1120_n_spl_
  );


  or

  (
    g1227_n,
    g1118_n_spl_,
    g1120_p_spl_
  );


  and

  (
    g1228_p,
    g1121_n_spl_,
    g1227_n
  );


  or

  (
    g1228_n,
    g1121_p_spl_,
    g1227_p
  );


  and

  (
    g1229_p,
    g1226_n_spl_,
    g1228_p_spl_
  );


  or

  (
    g1229_n,
    g1226_p_spl_,
    g1228_n_spl_
  );


  and

  (
    g1230_p,
    g1226_p_spl_,
    g1228_n_spl_
  );


  or

  (
    g1230_n,
    g1226_n_spl_,
    g1228_p_spl_
  );


  and

  (
    g1231_p,
    g1229_n_spl_,
    g1230_n
  );


  or

  (
    g1231_n,
    g1229_p_spl_,
    g1230_p
  );


  and

  (
    g1232_p,
    g1225_n_spl_,
    g1231_p_spl_
  );


  or

  (
    g1232_n,
    g1225_p_spl_,
    g1231_n_spl_
  );


  and

  (
    g1233_p,
    g1225_p_spl_,
    g1231_n_spl_
  );


  or

  (
    g1233_n,
    g1225_n_spl_,
    g1231_p_spl_
  );


  and

  (
    g1234_p,
    g1232_n_spl_,
    g1233_n
  );


  or

  (
    g1234_n,
    g1232_p_spl_,
    g1233_p
  );


  and

  (
    g1235_p,
    g1224_n_spl_,
    g1234_p_spl_
  );


  or

  (
    g1235_n,
    g1224_p_spl_,
    g1234_n_spl_
  );


  and

  (
    g1236_p,
    g1224_p_spl_,
    g1234_n_spl_
  );


  or

  (
    g1236_n,
    g1224_n_spl_,
    g1234_p_spl_
  );


  and

  (
    g1237_p,
    g1235_n_spl_,
    g1236_n
  );


  or

  (
    g1237_n,
    g1235_p_spl_,
    g1236_p
  );


  and

  (
    g1238_p,
    g1223_n_spl_,
    g1237_p_spl_
  );


  or

  (
    g1238_n,
    g1223_p_spl_,
    g1237_n_spl_
  );


  and

  (
    g1239_p,
    g1223_p_spl_,
    g1237_n_spl_
  );


  or

  (
    g1239_n,
    g1223_n_spl_,
    g1237_p_spl_
  );


  and

  (
    g1240_p,
    g1238_n_spl_,
    g1239_n
  );


  or

  (
    g1240_n,
    g1238_p_spl_,
    g1239_p
  );


  and

  (
    g1241_p,
    g1222_n_spl_,
    g1240_p_spl_
  );


  or

  (
    g1241_n,
    g1222_p_spl_,
    g1240_n_spl_
  );


  and

  (
    g1242_p,
    g988_n,
    g1012_p_spl_
  );


  or

  (
    g1242_n,
    g988_p_spl_,
    g1012_n
  );


  and

  (
    g1243_p,
    G3_p_spl_00,
    G17_p_spl_000
  );


  or

  (
    g1243_n,
    G3_n_spl_0,
    G17_n_spl_000
  );


  and

  (
    g1244_p,
    G2_p_spl_00,
    G18_p_spl_000
  );


  or

  (
    g1244_n,
    G2_n_spl_0,
    G18_n_spl_000
  );


  and

  (
    g1245_p,
    g1243_p_spl_,
    g1244_p_spl_
  );


  or

  (
    g1245_n,
    g1243_n_spl_,
    g1244_n_spl_
  );


  and

  (
    g1246_p,
    g1243_n_spl_,
    g1244_n_spl_
  );


  or

  (
    g1246_n,
    g1243_p_spl_,
    g1244_p_spl_
  );


  and

  (
    g1247_p,
    g1245_n_spl_0,
    g1246_n
  );


  or

  (
    g1247_n,
    g1245_p_spl_0,
    g1246_p
  );


  and

  (
    g1248_p,
    g989_n_spl_,
    g1247_n_spl_
  );


  or

  (
    g1248_n,
    g989_p_spl_0,
    g1247_p_spl_
  );


  and

  (
    g1249_p,
    g989_p_spl_0,
    g1247_p_spl_
  );


  or

  (
    g1249_n,
    g989_n_spl_,
    g1247_n_spl_
  );


  and

  (
    g1250_p,
    g1248_n_spl_,
    g1249_n
  );


  or

  (
    g1250_n,
    g1248_p_spl_,
    g1249_p
  );


  and

  (
    g1251_p,
    g982_n_spl_,
    g987_n
  );


  or

  (
    g1251_n,
    g982_p_spl_,
    g987_p_spl_
  );


  and

  (
    g1252_p,
    n2821_lo_p_spl_001,
    n6053_o2_p_spl_1
  );


  or

  (
    g1252_n,
    n2821_lo_n_spl_01,
    n6053_o2_n_spl_1
  );


  and

  (
    g1253_p,
    g976_n_spl_,
    g979_n_spl_
  );


  or

  (
    g1253_n,
    g976_p_spl_,
    g979_p_spl_
  );


  and

  (
    g1254_p,
    n2809_lo_p_spl_011,
    n6024_o2_p_spl_01
  );


  or

  (
    g1254_n,
    n2809_lo_n_spl_10,
    n6024_o2_n_spl_0
  );


  and

  (
    g1255_p,
    g970_n_spl_,
    g973_n_spl_
  );


  or

  (
    g1255_n,
    g970_p_spl_,
    g973_p_spl_
  );


  and

  (
    g1256_p,
    n2797_lo_p_spl_101,
    n6025_o2_p_spl_00
  );


  or

  (
    g1256_n,
    n2797_lo_n_spl_101,
    n6025_o2_n_spl_00
  );


  and

  (
    g1257_p,
    n1003_o2_p_spl_,
    g967_n_spl_
  );


  or

  (
    g1257_n,
    n1003_o2_n_spl_,
    g967_p_spl_
  );


  and

  (
    g1258_p,
    g1165_p_spl_,
    g1166_n_spl_
  );


  or

  (
    g1258_n,
    g1165_n_spl_,
    g1166_p_spl_
  );


  and

  (
    g1259_p,
    g1167_n_spl_,
    g1258_n
  );


  or

  (
    g1259_n,
    g1167_p_spl_,
    g1258_p
  );


  and

  (
    g1260_p,
    g1257_n_spl_,
    g1259_p_spl_
  );


  or

  (
    g1260_n,
    g1257_p_spl_,
    g1259_n_spl_
  );


  and

  (
    g1261_p,
    g1257_p_spl_,
    g1259_n_spl_
  );


  or

  (
    g1261_n,
    g1257_n_spl_,
    g1259_p_spl_
  );


  and

  (
    g1262_p,
    g1260_n_spl_,
    g1261_n
  );


  or

  (
    g1262_n,
    g1260_p_spl_,
    g1261_p
  );


  and

  (
    g1263_p,
    g1256_n_spl_,
    g1262_p_spl_
  );


  or

  (
    g1263_n,
    g1256_p_spl_,
    g1262_n_spl_
  );


  and

  (
    g1264_p,
    g1256_p_spl_,
    g1262_n_spl_
  );


  or

  (
    g1264_n,
    g1256_n_spl_,
    g1262_p_spl_
  );


  and

  (
    g1265_p,
    g1263_n_spl_,
    g1264_n
  );


  or

  (
    g1265_n,
    g1263_p_spl_,
    g1264_p
  );


  and

  (
    g1266_p,
    g1255_n_spl_,
    g1265_p_spl_
  );


  or

  (
    g1266_n,
    g1255_p_spl_,
    g1265_n_spl_
  );


  and

  (
    g1267_p,
    g1255_p_spl_,
    g1265_n_spl_
  );


  or

  (
    g1267_n,
    g1255_n_spl_,
    g1265_p_spl_
  );


  and

  (
    g1268_p,
    g1266_n_spl_,
    g1267_n
  );


  or

  (
    g1268_n,
    g1266_p_spl_,
    g1267_p
  );


  and

  (
    g1269_p,
    g1254_n_spl_,
    g1268_p_spl_
  );


  or

  (
    g1269_n,
    g1254_p_spl_,
    g1268_n_spl_
  );


  and

  (
    g1270_p,
    g1254_p_spl_,
    g1268_n_spl_
  );


  or

  (
    g1270_n,
    g1254_n_spl_,
    g1268_p_spl_
  );


  and

  (
    g1271_p,
    g1269_n_spl_,
    g1270_n
  );


  or

  (
    g1271_n,
    g1269_p_spl_,
    g1270_p
  );


  and

  (
    g1272_p,
    g1253_n_spl_,
    g1271_p_spl_
  );


  or

  (
    g1272_n,
    g1253_p_spl_,
    g1271_n_spl_
  );


  and

  (
    g1273_p,
    g1253_p_spl_,
    g1271_n_spl_
  );


  or

  (
    g1273_n,
    g1253_n_spl_,
    g1271_p_spl_
  );


  and

  (
    g1274_p,
    g1272_n_spl_,
    g1273_n
  );


  or

  (
    g1274_n,
    g1272_p_spl_,
    g1273_p
  );


  and

  (
    g1275_p,
    g1252_n_spl_,
    g1274_p_spl_
  );


  or

  (
    g1275_n,
    g1252_p_spl_,
    g1274_n_spl_
  );


  and

  (
    g1276_p,
    g1252_p_spl_,
    g1274_n_spl_
  );


  or

  (
    g1276_n,
    g1252_n_spl_,
    g1274_p_spl_
  );


  and

  (
    g1277_p,
    g1275_n_spl_,
    g1276_n
  );


  or

  (
    g1277_n,
    g1275_p_spl_,
    g1276_p
  );


  or

  (
    g1278_n,
    g1251_p,
    g1277_n
  );


  and

  (
    g1279_p,
    n1374_o2_n_spl_,
    n1392_o2_p_spl_
  );


  or

  (
    g1279_n,
    n1374_o2_p_spl_,
    n1392_o2_n_spl_
  );


  and

  (
    g1280_p,
    n1390_o2_p,
    g1279_n_spl_
  );


  or

  (
    g1280_n,
    n1390_o2_n,
    g1279_p_spl_
  );


  and

  (
    g1281_p,
    n1488_o2_n_spl_,
    n1501_o2_p_spl_
  );


  or

  (
    g1281_n,
    n1488_o2_p_spl_,
    n1501_o2_n_spl_
  );


  and

  (
    g1282_p,
    n1488_o2_p_spl_,
    n1501_o2_n_spl_
  );


  or

  (
    g1282_n,
    n1488_o2_n_spl_,
    n1501_o2_p_spl_
  );


  and

  (
    g1283_p,
    g1281_n_spl_,
    g1282_n
  );


  or

  (
    g1283_n,
    g1281_p_spl_,
    g1282_p
  );


  and

  (
    g1284_p,
    g1280_n_spl_,
    g1283_p_spl_
  );


  or

  (
    g1284_n,
    g1280_p_spl_,
    g1283_n_spl_
  );


  and

  (
    g1285_p,
    n2734_lo_p_spl_001,
    lo050_buf_o2_p_spl_0
  );


  or

  (
    g1285_n,
    n2734_lo_n_spl_001,
    lo050_buf_o2_n_spl_0
  );


  and

  (
    g1286_p,
    g1280_p_spl_,
    g1283_n_spl_
  );


  or

  (
    g1286_n,
    g1280_n_spl_,
    g1283_p_spl_
  );


  and

  (
    g1287_p,
    g1284_n_spl_,
    g1286_n
  );


  or

  (
    g1287_n,
    g1284_p_spl_,
    g1286_p
  );


  and

  (
    g1288_p,
    g1285_n_spl_,
    g1287_p_spl_
  );


  or

  (
    g1288_n,
    g1285_p_spl_,
    g1287_n_spl_
  );


  and

  (
    g1289_p,
    g1284_n_spl_,
    g1288_n_spl_
  );


  or

  (
    g1289_n,
    g1284_p_spl_,
    g1288_p_spl_
  );


  and

  (
    g1290_p,
    n2734_lo_p_spl_010,
    lo054_buf_o2_p_spl_0
  );


  or

  (
    g1290_n,
    n2734_lo_n_spl_010,
    lo054_buf_o2_n_spl_0
  );


  and

  (
    g1291_p,
    n1499_o2_p,
    g1281_n_spl_
  );


  or

  (
    g1291_n,
    n1499_o2_n,
    g1281_p_spl_
  );


  and

  (
    g1292_p,
    lo058_buf_o2_p_spl_0,
    lo082_buf_o2_p_spl_0
  );


  or

  (
    g1292_n,
    lo058_buf_o2_n_spl_0,
    lo082_buf_o2_n_spl_0
  );


  and

  (
    g1293_p,
    n1602_o2_n_spl_,
    n1603_o2_n_spl_
  );


  or

  (
    g1293_n,
    n1602_o2_p_spl_,
    n1603_o2_p_spl_
  );


  and

  (
    g1294_p,
    n1602_o2_p_spl_,
    n1603_o2_p_spl_
  );


  or

  (
    g1294_n,
    n1602_o2_n_spl_,
    n1603_o2_n_spl_
  );


  and

  (
    g1295_p,
    g1293_n_spl_,
    g1294_n
  );


  or

  (
    g1295_n,
    g1293_p_spl_,
    g1294_p
  );


  and

  (
    g1296_p,
    g1292_n_spl_,
    g1295_p_spl_
  );


  or

  (
    g1296_n,
    g1292_p_spl_,
    g1295_n_spl_
  );


  and

  (
    g1297_p,
    g1292_p_spl_,
    g1295_n_spl_
  );


  or

  (
    g1297_n,
    g1292_n_spl_,
    g1295_p_spl_
  );


  and

  (
    g1298_p,
    g1296_n_spl_,
    g1297_n
  );


  or

  (
    g1298_n,
    g1296_p_spl_,
    g1297_p
  );


  and

  (
    g1299_p,
    g1291_n_spl_,
    g1298_p_spl_
  );


  or

  (
    g1299_n,
    g1291_p_spl_,
    g1298_n_spl_
  );


  and

  (
    g1300_p,
    g1291_p_spl_,
    g1298_n_spl_
  );


  or

  (
    g1300_n,
    g1291_n_spl_,
    g1298_p_spl_
  );


  and

  (
    g1301_p,
    g1299_n_spl_,
    g1300_n
  );


  or

  (
    g1301_n,
    g1299_p_spl_,
    g1300_p
  );


  and

  (
    g1302_p,
    g1290_n_spl_,
    g1301_p_spl_
  );


  or

  (
    g1302_n,
    g1290_p_spl_,
    g1301_n_spl_
  );


  and

  (
    g1303_p,
    g1290_p_spl_,
    g1301_n_spl_
  );


  or

  (
    g1303_n,
    g1290_n_spl_,
    g1301_p_spl_
  );


  and

  (
    g1304_p,
    g1302_n_spl_,
    g1303_n
  );


  or

  (
    g1304_n,
    g1302_p_spl_,
    g1303_p
  );


  and

  (
    g1305_p,
    g1289_n_spl_,
    g1304_p_spl_
  );


  or

  (
    g1305_n,
    g1289_p_spl_,
    g1304_n_spl_
  );


  and

  (
    g1306_p,
    n2746_lo_p_spl_001,
    lo050_buf_o2_p_spl_0
  );


  or

  (
    g1306_n,
    n2746_lo_n_spl_001,
    lo050_buf_o2_n_spl_0
  );


  and

  (
    g1307_p,
    g1289_p_spl_,
    g1304_n_spl_
  );


  or

  (
    g1307_n,
    g1289_n_spl_,
    g1304_p_spl_
  );


  and

  (
    g1308_p,
    g1305_n_spl_,
    g1307_n
  );


  or

  (
    g1308_n,
    g1305_p_spl_,
    g1307_p
  );


  and

  (
    g1309_p,
    g1306_n_spl_,
    g1308_p_spl_
  );


  or

  (
    g1309_n,
    g1306_p_spl_,
    g1308_n_spl_
  );


  and

  (
    g1310_p,
    g1305_n_spl_,
    g1309_n_spl_
  );


  or

  (
    g1310_n,
    g1305_p_spl_,
    g1309_p_spl_
  );


  and

  (
    g1311_p,
    n2746_lo_p_spl_001,
    lo054_buf_o2_p_spl_0
  );


  or

  (
    g1311_n,
    n2746_lo_n_spl_001,
    lo054_buf_o2_n_spl_0
  );


  and

  (
    g1312_p,
    g1299_n_spl_,
    g1302_n_spl_
  );


  or

  (
    g1312_n,
    g1299_p_spl_,
    g1302_p_spl_
  );


  and

  (
    g1313_p,
    n2734_lo_p_spl_010,
    lo058_buf_o2_p_spl_0
  );


  or

  (
    g1313_n,
    n2734_lo_n_spl_010,
    lo058_buf_o2_n_spl_0
  );


  and

  (
    g1314_p,
    lo062_buf_o2_p_spl_0,
    lo082_buf_o2_p_spl_
  );


  or

  (
    g1314_n,
    lo062_buf_o2_n_spl_0,
    lo082_buf_o2_n_spl_
  );


  and

  (
    g1315_p,
    g1293_n_spl_,
    g1296_n_spl_
  );


  or

  (
    g1315_n,
    g1293_p_spl_,
    g1296_p_spl_
  );


  and

  (
    g1316_p,
    g1314_n_spl_,
    g1315_n_spl_
  );


  or

  (
    g1316_n,
    g1314_p_spl_,
    g1315_p_spl_
  );


  and

  (
    g1317_p,
    g1314_p_spl_,
    g1315_p_spl_
  );


  or

  (
    g1317_n,
    g1314_n_spl_,
    g1315_n_spl_
  );


  and

  (
    g1318_p,
    g1316_n_spl_,
    g1317_n
  );


  or

  (
    g1318_n,
    g1316_p_spl_,
    g1317_p
  );


  and

  (
    g1319_p,
    g1313_n_spl_,
    g1318_p_spl_
  );


  or

  (
    g1319_n,
    g1313_p_spl_,
    g1318_n_spl_
  );


  and

  (
    g1320_p,
    g1313_p_spl_,
    g1318_n_spl_
  );


  or

  (
    g1320_n,
    g1313_n_spl_,
    g1318_p_spl_
  );


  and

  (
    g1321_p,
    g1319_n_spl_,
    g1320_n
  );


  or

  (
    g1321_n,
    g1319_p_spl_,
    g1320_p
  );


  and

  (
    g1322_p,
    g1312_n_spl_,
    g1321_p_spl_
  );


  or

  (
    g1322_n,
    g1312_p_spl_,
    g1321_n_spl_
  );


  and

  (
    g1323_p,
    g1312_p_spl_,
    g1321_n_spl_
  );


  or

  (
    g1323_n,
    g1312_n_spl_,
    g1321_p_spl_
  );


  and

  (
    g1324_p,
    g1322_n_spl_,
    g1323_n
  );


  or

  (
    g1324_n,
    g1322_p_spl_,
    g1323_p
  );


  and

  (
    g1325_p,
    g1311_n_spl_,
    g1324_p_spl_
  );


  or

  (
    g1325_n,
    g1311_p_spl_,
    g1324_n_spl_
  );


  and

  (
    g1326_p,
    g1311_p_spl_,
    g1324_n_spl_
  );


  or

  (
    g1326_n,
    g1311_n_spl_,
    g1324_p_spl_
  );


  and

  (
    g1327_p,
    g1325_n_spl_,
    g1326_n
  );


  or

  (
    g1327_n,
    g1325_p_spl_,
    g1326_p
  );


  and

  (
    g1328_p,
    g1310_n_spl_,
    g1327_p_spl_
  );


  or

  (
    g1328_n,
    g1310_p_spl_,
    g1327_n_spl_
  );


  and

  (
    g1329_p,
    n1045_o2_n_spl_,
    n1069_o2_p_spl_
  );


  or

  (
    g1329_n,
    n1045_o2_p_spl_,
    n1069_o2_n_spl_
  );


  and

  (
    g1330_p,
    n1067_o2_p,
    g1329_n_spl_
  );


  or

  (
    g1330_n,
    n1067_o2_n,
    g1329_p_spl_
  );


  and

  (
    g1331_p,
    n1147_o2_n_spl_,
    n1171_o2_p_spl_
  );


  or

  (
    g1331_n,
    n1147_o2_p_spl_,
    n1171_o2_n_spl_
  );


  and

  (
    g1332_p,
    n1147_o2_p_spl_,
    n1171_o2_n_spl_
  );


  or

  (
    g1332_n,
    n1147_o2_n_spl_,
    n1171_o2_p_spl_
  );


  and

  (
    g1333_p,
    g1331_n_spl_,
    g1332_n
  );


  or

  (
    g1333_n,
    g1331_p_spl_,
    g1332_p
  );


  and

  (
    g1334_p,
    g1330_n_spl_,
    g1333_p_spl_
  );


  or

  (
    g1334_n,
    g1330_p_spl_,
    g1333_n_spl_
  );


  and

  (
    g1335_p,
    n2734_lo_p_spl_011,
    lo038_buf_o2_p_spl_00
  );


  or

  (
    g1335_n,
    n2734_lo_n_spl_011,
    lo038_buf_o2_n_spl_0
  );


  and

  (
    g1336_p,
    g1330_p_spl_,
    g1333_n_spl_
  );


  or

  (
    g1336_n,
    g1330_n_spl_,
    g1333_p_spl_
  );


  and

  (
    g1337_p,
    g1334_n_spl_,
    g1336_n
  );


  or

  (
    g1337_n,
    g1334_p_spl_,
    g1336_p
  );


  and

  (
    g1338_p,
    g1335_n_spl_,
    g1337_p_spl_
  );


  or

  (
    g1338_n,
    g1335_p_spl_,
    g1337_n_spl_
  );


  and

  (
    g1339_p,
    g1334_n_spl_,
    g1338_n_spl_
  );


  or

  (
    g1339_n,
    g1334_p_spl_,
    g1338_p_spl_
  );


  and

  (
    g1340_p,
    n2734_lo_p_spl_011,
    lo042_buf_o2_p_spl_0
  );


  or

  (
    g1340_n,
    n2734_lo_n_spl_011,
    lo042_buf_o2_n_spl_0
  );


  and

  (
    g1341_p,
    n1169_o2_p,
    g1331_n_spl_
  );


  or

  (
    g1341_n,
    n1169_o2_n,
    g1331_p_spl_
  );


  and

  (
    g1342_p,
    n1257_o2_n_spl_,
    n1281_o2_p_spl_
  );


  or

  (
    g1342_n,
    n1257_o2_p_spl_,
    n1281_o2_n_spl_
  );


  and

  (
    g1343_p,
    n1257_o2_p_spl_,
    n1281_o2_n_spl_
  );


  or

  (
    g1343_n,
    n1257_o2_n_spl_,
    n1281_o2_p_spl_
  );


  and

  (
    g1344_p,
    g1342_n_spl_,
    g1343_n
  );


  or

  (
    g1344_n,
    g1342_p_spl_,
    g1343_p
  );


  and

  (
    g1345_p,
    g1341_n_spl_,
    g1344_p_spl_
  );


  or

  (
    g1345_n,
    g1341_p_spl_,
    g1344_n_spl_
  );


  and

  (
    g1346_p,
    g1341_p_spl_,
    g1344_n_spl_
  );


  or

  (
    g1346_n,
    g1341_n_spl_,
    g1344_p_spl_
  );


  and

  (
    g1347_p,
    g1345_n_spl_,
    g1346_n
  );


  or

  (
    g1347_n,
    g1345_p_spl_,
    g1346_p
  );


  and

  (
    g1348_p,
    g1340_n_spl_,
    g1347_p_spl_
  );


  or

  (
    g1348_n,
    g1340_p_spl_,
    g1347_n_spl_
  );


  and

  (
    g1349_p,
    g1340_p_spl_,
    g1347_n_spl_
  );


  or

  (
    g1349_n,
    g1340_n_spl_,
    g1347_p_spl_
  );


  and

  (
    g1350_p,
    g1348_n_spl_,
    g1349_n
  );


  or

  (
    g1350_n,
    g1348_p_spl_,
    g1349_p
  );


  and

  (
    g1351_p,
    g1339_n_spl_,
    g1350_p_spl_
  );


  or

  (
    g1351_n,
    g1339_p_spl_,
    g1350_n_spl_
  );


  and

  (
    g1352_p,
    n2746_lo_p_spl_010,
    lo038_buf_o2_p_spl_00
  );


  or

  (
    g1352_n,
    n2746_lo_n_spl_010,
    lo038_buf_o2_n_spl_0
  );


  and

  (
    g1353_p,
    g1339_p_spl_,
    g1350_n_spl_
  );


  or

  (
    g1353_n,
    g1339_n_spl_,
    g1350_p_spl_
  );


  and

  (
    g1354_p,
    g1351_n_spl_,
    g1353_n
  );


  or

  (
    g1354_n,
    g1351_p_spl_,
    g1353_p
  );


  and

  (
    g1355_p,
    g1352_n_spl_,
    g1354_p_spl_
  );


  or

  (
    g1355_n,
    g1352_p_spl_,
    g1354_n_spl_
  );


  and

  (
    g1356_p,
    g1351_n_spl_,
    g1355_n_spl_
  );


  or

  (
    g1356_n,
    g1351_p_spl_,
    g1355_p_spl_
  );


  and

  (
    g1357_p,
    n2746_lo_p_spl_010,
    lo042_buf_o2_p_spl_0
  );


  or

  (
    g1357_n,
    n2746_lo_n_spl_010,
    lo042_buf_o2_n_spl_0
  );


  and

  (
    g1358_p,
    g1345_n_spl_,
    g1348_n_spl_
  );


  or

  (
    g1358_n,
    g1345_p_spl_,
    g1348_p_spl_
  );


  and

  (
    g1359_p,
    n2734_lo_p_spl_100,
    lo046_buf_o2_p_spl_0
  );


  or

  (
    g1359_n,
    n2734_lo_n_spl_100,
    lo046_buf_o2_n_spl_0
  );


  and

  (
    g1360_p,
    n1279_o2_p,
    g1342_n_spl_
  );


  or

  (
    g1360_n,
    n1279_o2_n,
    g1342_p_spl_
  );


  and

  (
    g1361_p,
    n1374_o2_p_spl_,
    n1392_o2_n_spl_
  );


  or

  (
    g1361_n,
    n1374_o2_n_spl_,
    n1392_o2_p_spl_
  );


  and

  (
    g1362_p,
    g1279_n_spl_,
    g1361_n
  );


  or

  (
    g1362_n,
    g1279_p_spl_,
    g1361_p
  );


  and

  (
    g1363_p,
    g1360_n_spl_,
    g1362_p_spl_
  );


  or

  (
    g1363_n,
    g1360_p_spl_,
    g1362_n_spl_
  );


  and

  (
    g1364_p,
    g1360_p_spl_,
    g1362_n_spl_
  );


  or

  (
    g1364_n,
    g1360_n_spl_,
    g1362_p_spl_
  );


  and

  (
    g1365_p,
    g1363_n_spl_,
    g1364_n
  );


  or

  (
    g1365_n,
    g1363_p_spl_,
    g1364_p
  );


  and

  (
    g1366_p,
    g1359_n_spl_,
    g1365_p_spl_
  );


  or

  (
    g1366_n,
    g1359_p_spl_,
    g1365_n_spl_
  );


  and

  (
    g1367_p,
    g1359_p_spl_,
    g1365_n_spl_
  );


  or

  (
    g1367_n,
    g1359_n_spl_,
    g1365_p_spl_
  );


  and

  (
    g1368_p,
    g1366_n_spl_,
    g1367_n
  );


  or

  (
    g1368_n,
    g1366_p_spl_,
    g1367_p
  );


  and

  (
    g1369_p,
    g1358_n_spl_,
    g1368_p_spl_
  );


  or

  (
    g1369_n,
    g1358_p_spl_,
    g1368_n_spl_
  );


  and

  (
    g1370_p,
    g1358_p_spl_,
    g1368_n_spl_
  );


  or

  (
    g1370_n,
    g1358_n_spl_,
    g1368_p_spl_
  );


  and

  (
    g1371_p,
    g1369_n_spl_,
    g1370_n
  );


  or

  (
    g1371_n,
    g1369_p_spl_,
    g1370_p
  );


  and

  (
    g1372_p,
    g1357_n_spl_,
    g1371_p_spl_
  );


  or

  (
    g1372_n,
    g1357_p_spl_,
    g1371_n_spl_
  );


  and

  (
    g1373_p,
    g1357_p_spl_,
    g1371_n_spl_
  );


  or

  (
    g1373_n,
    g1357_n_spl_,
    g1371_p_spl_
  );


  and

  (
    g1374_p,
    g1372_n_spl_,
    g1373_n
  );


  or

  (
    g1374_n,
    g1372_p_spl_,
    g1373_p
  );


  and

  (
    g1375_p,
    g1356_n_spl_,
    g1374_p_spl_
  );


  or

  (
    g1375_n,
    g1356_p_spl_,
    g1374_n_spl_
  );


  and

  (
    g1376_p,
    n2758_lo_p_spl_000,
    lo038_buf_o2_p_spl_0
  );


  or

  (
    g1376_n,
    n2758_lo_n_spl_000,
    lo038_buf_o2_n_spl_1
  );


  and

  (
    g1377_p,
    g1356_p_spl_,
    g1374_n_spl_
  );


  or

  (
    g1377_n,
    g1356_n_spl_,
    g1374_p_spl_
  );


  and

  (
    g1378_p,
    g1375_n_spl_,
    g1377_n
  );


  or

  (
    g1378_n,
    g1375_p_spl_,
    g1377_p
  );


  and

  (
    g1379_p,
    g1376_n_spl_,
    g1378_p_spl_
  );


  or

  (
    g1379_n,
    g1376_p_spl_,
    g1378_n_spl_
  );


  and

  (
    g1380_p,
    g1375_n_spl_,
    g1379_n_spl_
  );


  or

  (
    g1380_n,
    g1375_p_spl_,
    g1379_p_spl_
  );


  and

  (
    g1381_p,
    n2758_lo_p_spl_001,
    lo042_buf_o2_p_spl_1
  );


  or

  (
    g1381_n,
    n2758_lo_n_spl_001,
    lo042_buf_o2_n_spl_1
  );


  and

  (
    g1382_p,
    g1369_n_spl_,
    g1372_n_spl_
  );


  or

  (
    g1382_n,
    g1369_p_spl_,
    g1372_p_spl_
  );


  and

  (
    g1383_p,
    n2746_lo_p_spl_011,
    lo046_buf_o2_p_spl_0
  );


  or

  (
    g1383_n,
    n2746_lo_n_spl_011,
    lo046_buf_o2_n_spl_0
  );


  and

  (
    g1384_p,
    g1363_n_spl_,
    g1366_n_spl_
  );


  or

  (
    g1384_n,
    g1363_p_spl_,
    g1366_p_spl_
  );


  and

  (
    g1385_p,
    g1285_p_spl_,
    g1287_n_spl_
  );


  or

  (
    g1385_n,
    g1285_n_spl_,
    g1287_p_spl_
  );


  and

  (
    g1386_p,
    g1288_n_spl_,
    g1385_n
  );


  or

  (
    g1386_n,
    g1288_p_spl_,
    g1385_p
  );


  and

  (
    g1387_p,
    g1384_n_spl_,
    g1386_p_spl_
  );


  or

  (
    g1387_n,
    g1384_p_spl_,
    g1386_n_spl_
  );


  and

  (
    g1388_p,
    g1384_p_spl_,
    g1386_n_spl_
  );


  or

  (
    g1388_n,
    g1384_n_spl_,
    g1386_p_spl_
  );


  and

  (
    g1389_p,
    g1387_n_spl_,
    g1388_n
  );


  or

  (
    g1389_n,
    g1387_p_spl_,
    g1388_p
  );


  and

  (
    g1390_p,
    g1383_n_spl_,
    g1389_p_spl_
  );


  or

  (
    g1390_n,
    g1383_p_spl_,
    g1389_n_spl_
  );


  and

  (
    g1391_p,
    g1383_p_spl_,
    g1389_n_spl_
  );


  or

  (
    g1391_n,
    g1383_n_spl_,
    g1389_p_spl_
  );


  and

  (
    g1392_p,
    g1390_n_spl_,
    g1391_n
  );


  or

  (
    g1392_n,
    g1390_p_spl_,
    g1391_p
  );


  and

  (
    g1393_p,
    g1382_n_spl_,
    g1392_p_spl_
  );


  or

  (
    g1393_n,
    g1382_p_spl_,
    g1392_n_spl_
  );


  and

  (
    g1394_p,
    g1382_p_spl_,
    g1392_n_spl_
  );


  or

  (
    g1394_n,
    g1382_n_spl_,
    g1392_p_spl_
  );


  and

  (
    g1395_p,
    g1393_n_spl_,
    g1394_n
  );


  or

  (
    g1395_n,
    g1393_p_spl_,
    g1394_p
  );


  and

  (
    g1396_p,
    g1381_n_spl_,
    g1395_p_spl_
  );


  or

  (
    g1396_n,
    g1381_p_spl_,
    g1395_n_spl_
  );


  and

  (
    g1397_p,
    g1381_p_spl_,
    g1395_n_spl_
  );


  or

  (
    g1397_n,
    g1381_n_spl_,
    g1395_p_spl_
  );


  and

  (
    g1398_p,
    g1396_n_spl_,
    g1397_n
  );


  or

  (
    g1398_n,
    g1396_p_spl_,
    g1397_p
  );


  and

  (
    g1399_p,
    g1380_n_spl_,
    g1398_p_spl_
  );


  or

  (
    g1399_n,
    g1380_p_spl_,
    g1398_n_spl_
  );


  and

  (
    g1400_p,
    g1016_n,
    g1250_p_spl_
  );


  or

  (
    g1400_n,
    g1016_p_spl_,
    g1250_n
  );


  or

  (
    g1401_n,
    n2833_lo_n_spl_00,
    n6148_o2_n_spl_1
  );


  or

  (
    g1402_n,
    n2770_lo_n_spl_000,
    lo002_buf_o2_n_spl_1
  );


  or

  (
    g1403_n,
    G1_n_spl_,
    G20_n_spl_000
  );


  or

  (
    g1404_n,
    n2860_lo_n_spl_11,
    n4842_o2_n_spl_
  );


  or

  (
    g1405_n,
    g935_n,
    g945_p
  );


  and

  (
    g1406_p,
    g946_n_spl_,
    g1405_n
  );


  and

  (
    g1407_p,
    g1404_n_spl_,
    g1406_p_spl_
  );


  or

  (
    g1408_n,
    g1404_n_spl_,
    g1406_p_spl_
  );


  or

  (
    g1409_n,
    n2848_lo_n_spl_11,
    n4845_o2_n_spl_
  );


  or

  (
    g1410_n,
    g923_n,
    g933_p
  );


  and

  (
    g1411_p,
    g934_n_spl_,
    g1410_n
  );


  and

  (
    g1412_p,
    g1409_n_spl_,
    g1411_p_spl_
  );


  or

  (
    g1413_n,
    g1409_n_spl_,
    g1411_p_spl_
  );


  or

  (
    g1414_n,
    n4848_o2_n_spl_,
    lo118_buf_o2_n_spl_11
  );


  or

  (
    g1415_n,
    g920_n,
    g921_n
  );


  and

  (
    g1416_p,
    g922_n_spl_,
    g1415_n
  );


  and

  (
    g1417_p,
    g1414_n_spl_,
    g1416_p_spl_
  );


  or

  (
    g1418_n,
    g1414_n_spl_,
    g1416_p_spl_
  );


  or

  (
    g1419_n,
    g928_p_spl_,
    g931_p_spl_
  );


  or

  (
    g1420_n,
    g916_n,
    g918_p
  );


  and

  (
    g1421_p,
    g919_n_spl_,
    g1420_n
  );


  and

  (
    g1422_p,
    g1419_n_spl_,
    g1421_p_spl_
  );


  or

  (
    g1423_n,
    g1419_n_spl_,
    g1421_p_spl_
  );


  or

  (
    g1424_n,
    g940_p_spl_,
    g943_p_spl_
  );


  or

  (
    g1425_n,
    g912_n,
    g914_p
  );


  and

  (
    g1426_p,
    g915_n_spl_,
    g1425_n
  );


  and

  (
    g1427_p,
    g1424_n_spl_,
    g1426_p_spl_
  );


  or

  (
    g1428_n,
    g1424_n_spl_,
    g1426_p_spl_
  );


  or

  (
    g1429_n,
    g952_p_spl_,
    g955_p_spl_
  );


  or

  (
    g1430_n,
    g908_n,
    g910_p
  );


  and

  (
    g1431_p,
    g911_n_spl_,
    g1430_n
  );


  and

  (
    g1432_p,
    g1429_n_spl_,
    g1431_p_spl_
  );


  or

  (
    g1433_n,
    g1429_n_spl_,
    g1431_p_spl_
  );


  and

  (
    g1434_p,
    g1013_n_spl_,
    g1015_p_spl_
  );


  and

  (
    g1435_p,
    n2833_lo_p_spl_00,
    n6026_o2_p_spl_1
  );


  or

  (
    g1435_n,
    n2833_lo_n_spl_00,
    n6026_o2_n_spl_1
  );


  and

  (
    g1436_p,
    g1222_p_spl_,
    g1240_n_spl_
  );


  or

  (
    g1436_n,
    g1222_n_spl_,
    g1240_p_spl_
  );


  and

  (
    g1437_p,
    g1241_n_spl_,
    g1436_n
  );


  or

  (
    g1437_n,
    g1241_p,
    g1436_p
  );


  or

  (
    g1438_n,
    g1435_p,
    g1437_n
  );


  and

  (
    g1439_p,
    n2821_lo_p_spl_01,
    n6029_o2_p_spl_1
  );


  or

  (
    g1439_n,
    n2821_lo_n_spl_10,
    n6029_o2_n_spl_1
  );


  and

  (
    g1440_p,
    g1145_p_spl_,
    g1163_n_spl_
  );


  or

  (
    g1440_n,
    g1145_n_spl_,
    g1163_p_spl_
  );


  and

  (
    g1441_p,
    g1164_n_spl_,
    g1440_n
  );


  or

  (
    g1441_n,
    g1164_p,
    g1440_p
  );


  or

  (
    g1442_n,
    g1439_p,
    g1441_n
  );


  and

  (
    g1443_p,
    n2809_lo_p_spl_100,
    n6032_o2_p_spl_1
  );


  or

  (
    g1443_n,
    n2809_lo_n_spl_10,
    n6032_o2_n_spl_
  );


  and

  (
    g1444_p,
    g1088_p_spl_,
    g1106_n_spl_
  );


  or

  (
    g1444_n,
    g1088_n_spl_,
    g1106_p_spl_
  );


  and

  (
    g1445_p,
    g1107_n_spl_,
    g1444_n
  );


  or

  (
    g1445_n,
    g1107_p,
    g1444_p
  );


  or

  (
    g1446_n,
    g1443_p,
    g1445_n
  );


  and

  (
    g1447_p,
    n2797_lo_p_spl_110,
    n6035_o2_p_spl_1
  );


  or

  (
    g1447_n,
    n2797_lo_n_spl_11,
    n6035_o2_n_spl_
  );


  and

  (
    g1448_p,
    g1043_p_spl_,
    g1052_n_spl_
  );


  or

  (
    g1448_n,
    g1043_n_spl_,
    g1052_p_spl_
  );


  and

  (
    g1449_p,
    g1053_n_spl_,
    g1448_n
  );


  or

  (
    g1449_n,
    g1053_p,
    g1448_p
  );


  or

  (
    g1450_n,
    g1447_p,
    g1449_n
  );


  and

  (
    g1451_p,
    n6037_o2_p_spl_1,
    lo102_buf_o2_p_spl_111
  );


  or

  (
    g1451_n,
    n6037_o2_n_spl_,
    lo102_buf_o2_n_spl_111
  );


  and

  (
    g1452_p,
    g1047_n_spl_,
    g1050_n_spl_
  );


  or

  (
    g1452_n,
    g1047_p_spl_,
    g1050_p_spl_
  );


  or

  (
    g1453_n,
    g1451_p,
    g1452_p
  );


  or

  (
    g1454_n,
    n2833_lo_n_spl_0,
    n6053_o2_n_spl_1
  );


  and

  (
    g1455_p,
    g1272_n_spl_,
    g1275_n_spl_
  );


  or

  (
    g1455_n,
    g1272_p_spl_,
    g1275_p_spl_
  );


  and

  (
    g1456_p,
    n2821_lo_p_spl_01,
    n6024_o2_p_spl_01
  );


  or

  (
    g1456_n,
    n2821_lo_n_spl_10,
    n6024_o2_n_spl_1
  );


  and

  (
    g1457_p,
    g1266_n_spl_,
    g1269_n_spl_
  );


  or

  (
    g1457_n,
    g1266_p_spl_,
    g1269_p_spl_
  );


  and

  (
    g1458_p,
    n2809_lo_p_spl_100,
    n6025_o2_p_spl_01
  );


  or

  (
    g1458_n,
    n2809_lo_n_spl_11,
    n6025_o2_n_spl_0
  );


  and

  (
    g1459_p,
    g1260_n_spl_,
    g1263_n_spl_
  );


  or

  (
    g1459_n,
    g1260_p_spl_,
    g1263_p_spl_
  );


  and

  (
    g1460_p,
    g1175_p_spl_,
    g1177_n_spl_
  );


  or

  (
    g1460_n,
    g1175_n_spl_,
    g1177_p_spl_
  );


  and

  (
    g1461_p,
    g1178_n_spl_,
    g1460_n
  );


  or

  (
    g1461_n,
    g1178_p_spl_,
    g1460_p
  );


  and

  (
    g1462_p,
    g1459_n_spl_,
    g1461_p_spl_
  );


  or

  (
    g1462_n,
    g1459_p_spl_,
    g1461_n_spl_
  );


  and

  (
    g1463_p,
    g1459_p_spl_,
    g1461_n_spl_
  );


  or

  (
    g1463_n,
    g1459_n_spl_,
    g1461_p_spl_
  );


  and

  (
    g1464_p,
    g1462_n_spl_,
    g1463_n
  );


  or

  (
    g1464_n,
    g1462_p_spl_,
    g1463_p
  );


  and

  (
    g1465_p,
    g1458_n_spl_,
    g1464_p_spl_
  );


  or

  (
    g1465_n,
    g1458_p_spl_,
    g1464_n_spl_
  );


  and

  (
    g1466_p,
    g1458_p_spl_,
    g1464_n_spl_
  );


  or

  (
    g1466_n,
    g1458_n_spl_,
    g1464_p_spl_
  );


  and

  (
    g1467_p,
    g1465_n_spl_,
    g1466_n
  );


  or

  (
    g1467_n,
    g1465_p_spl_,
    g1466_p
  );


  and

  (
    g1468_p,
    g1457_n_spl_,
    g1467_p_spl_
  );


  or

  (
    g1468_n,
    g1457_p_spl_,
    g1467_n_spl_
  );


  and

  (
    g1469_p,
    g1457_p_spl_,
    g1467_n_spl_
  );


  or

  (
    g1469_n,
    g1457_n_spl_,
    g1467_p_spl_
  );


  and

  (
    g1470_p,
    g1468_n_spl_,
    g1469_n
  );


  or

  (
    g1470_n,
    g1468_p_spl_,
    g1469_p
  );


  and

  (
    g1471_p,
    g1456_n_spl_,
    g1470_p_spl_
  );


  or

  (
    g1471_n,
    g1456_p_spl_,
    g1470_n_spl_
  );


  and

  (
    g1472_p,
    g1456_p_spl_,
    g1470_n_spl_
  );


  or

  (
    g1472_n,
    g1456_n_spl_,
    g1470_p_spl_
  );


  and

  (
    g1473_p,
    g1471_n_spl_,
    g1472_n
  );


  or

  (
    g1473_n,
    g1471_p_spl_,
    g1472_p
  );


  and

  (
    g1474_p,
    g1455_n_spl_,
    g1473_p_spl_
  );


  or

  (
    g1474_n,
    g1455_p,
    g1473_n
  );


  or

  (
    g1475_n,
    g1455_n_spl_,
    g1473_p_spl_
  );


  and

  (
    g1476_p,
    g1474_n,
    g1475_n
  );


  and

  (
    g1477_p,
    g1454_n_spl_,
    g1476_p_spl_
  );


  and

  (
    g1478_p,
    g1101_n_spl_,
    g1104_n_spl_
  );


  or

  (
    g1478_n,
    g1101_p_spl_,
    g1104_p_spl_
  );


  and

  (
    g1479_p,
    n2797_lo_p_spl_110,
    n6034_o2_p_spl_1
  );


  or

  (
    g1479_n,
    n2797_lo_n_spl_11,
    n6034_o2_n_spl_
  );


  and

  (
    g1480_p,
    g1095_n_spl_,
    g1098_n_spl_
  );


  or

  (
    g1480_n,
    g1095_p_spl_,
    g1098_p_spl_
  );


  and

  (
    g1481_p,
    g1039_p_spl_,
    g1041_n_spl_
  );


  or

  (
    g1481_n,
    g1039_n_spl_,
    g1041_p_spl_
  );


  and

  (
    g1482_p,
    g1042_n_spl_,
    g1481_n
  );


  or

  (
    g1482_n,
    g1042_p_spl_,
    g1481_p
  );


  and

  (
    g1483_p,
    g1480_n_spl_,
    g1482_p_spl_
  );


  or

  (
    g1483_n,
    g1480_p_spl_,
    g1482_n_spl_
  );


  and

  (
    g1484_p,
    g1480_p_spl_,
    g1482_n_spl_
  );


  or

  (
    g1484_n,
    g1480_n_spl_,
    g1482_p_spl_
  );


  and

  (
    g1485_p,
    g1483_n_spl_,
    g1484_n
  );


  or

  (
    g1485_n,
    g1483_p,
    g1484_p
  );


  and

  (
    g1486_p,
    g1479_n_spl_,
    g1485_p_spl_
  );


  or

  (
    g1486_n,
    g1479_p_spl_,
    g1485_n_spl_
  );


  and

  (
    g1487_p,
    g1479_p_spl_,
    g1485_n_spl_
  );


  or

  (
    g1487_n,
    g1479_n_spl_,
    g1485_p_spl_
  );


  and

  (
    g1488_p,
    g1486_n_spl_,
    g1487_n
  );


  or

  (
    g1488_n,
    g1486_p,
    g1487_p
  );


  or

  (
    g1489_n,
    g1478_p,
    g1488_n
  );


  and

  (
    g1490_p,
    g1158_n_spl_,
    g1161_n_spl_
  );


  or

  (
    g1490_n,
    g1158_p_spl_,
    g1161_p_spl_
  );


  and

  (
    g1491_p,
    n2809_lo_p_spl_10,
    n6031_o2_p_spl_1
  );


  or

  (
    g1491_n,
    n2809_lo_n_spl_11,
    n6031_o2_n_spl_
  );


  and

  (
    g1492_p,
    g1152_n_spl_,
    g1155_n_spl_
  );


  or

  (
    g1492_n,
    g1152_p_spl_,
    g1155_p_spl_
  );


  and

  (
    g1493_p,
    g1084_p_spl_,
    g1086_n_spl_
  );


  or

  (
    g1493_n,
    g1084_n_spl_,
    g1086_p_spl_
  );


  and

  (
    g1494_p,
    g1087_n_spl_,
    g1493_n
  );


  or

  (
    g1494_n,
    g1087_p_spl_,
    g1493_p
  );


  and

  (
    g1495_p,
    g1492_n_spl_,
    g1494_p_spl_
  );


  or

  (
    g1495_n,
    g1492_p_spl_,
    g1494_n_spl_
  );


  and

  (
    g1496_p,
    g1492_p_spl_,
    g1494_n_spl_
  );


  or

  (
    g1496_n,
    g1492_n_spl_,
    g1494_p_spl_
  );


  and

  (
    g1497_p,
    g1495_n_spl_,
    g1496_n
  );


  or

  (
    g1497_n,
    g1495_p,
    g1496_p
  );


  and

  (
    g1498_p,
    g1491_n_spl_,
    g1497_p_spl_
  );


  or

  (
    g1498_n,
    g1491_p_spl_,
    g1497_n_spl_
  );


  and

  (
    g1499_p,
    g1491_p_spl_,
    g1497_n_spl_
  );


  or

  (
    g1499_n,
    g1491_n_spl_,
    g1497_p_spl_
  );


  and

  (
    g1500_p,
    g1498_n_spl_,
    g1499_n
  );


  or

  (
    g1500_n,
    g1498_p,
    g1499_p
  );


  or

  (
    g1501_n,
    g1490_p,
    g1500_n
  );


  and

  (
    g1502_p,
    g1235_n_spl_,
    g1238_n_spl_
  );


  or

  (
    g1502_n,
    g1235_p_spl_,
    g1238_p_spl_
  );


  and

  (
    g1503_p,
    n2821_lo_p_spl_10,
    n6028_o2_p_spl_1
  );


  or

  (
    g1503_n,
    n2821_lo_n_spl_11,
    n6028_o2_n_spl_1
  );


  and

  (
    g1504_p,
    g1229_n_spl_,
    g1232_n_spl_
  );


  or

  (
    g1504_n,
    g1229_p_spl_,
    g1232_p_spl_
  );


  and

  (
    g1505_p,
    g1141_p_spl_,
    g1143_n_spl_
  );


  or

  (
    g1505_n,
    g1141_n_spl_,
    g1143_p_spl_
  );


  and

  (
    g1506_p,
    g1144_n_spl_,
    g1505_n
  );


  or

  (
    g1506_n,
    g1144_p_spl_,
    g1505_p
  );


  and

  (
    g1507_p,
    g1504_n_spl_,
    g1506_p_spl_
  );


  or

  (
    g1507_n,
    g1504_p_spl_,
    g1506_n_spl_
  );


  and

  (
    g1508_p,
    g1504_p_spl_,
    g1506_n_spl_
  );


  or

  (
    g1508_n,
    g1504_n_spl_,
    g1506_p_spl_
  );


  and

  (
    g1509_p,
    g1507_n_spl_,
    g1508_n
  );


  or

  (
    g1509_n,
    g1507_p,
    g1508_p
  );


  and

  (
    g1510_p,
    g1503_n_spl_,
    g1509_p_spl_
  );


  or

  (
    g1510_n,
    g1503_p_spl_,
    g1509_n_spl_
  );


  and

  (
    g1511_p,
    g1503_p_spl_,
    g1509_n_spl_
  );


  or

  (
    g1511_n,
    g1503_n_spl_,
    g1509_p_spl_
  );


  and

  (
    g1512_p,
    g1510_n_spl_,
    g1511_n
  );


  or

  (
    g1512_n,
    g1510_p,
    g1511_p
  );


  or

  (
    g1513_n,
    g1502_p,
    g1512_n
  );


  or

  (
    g1514_n,
    g1251_n,
    g1277_p
  );


  and

  (
    g1515_p,
    g1278_n_spl_,
    g1514_n
  );


  and

  (
    g1516_p,
    n2770_lo_p_spl_000,
    lo038_buf_o2_p_spl_1
  );


  or

  (
    g1516_n,
    n2770_lo_n_spl_000,
    lo038_buf_o2_n_spl_1
  );


  and

  (
    g1517_p,
    g1380_p_spl_,
    g1398_n_spl_
  );


  or

  (
    g1517_n,
    g1380_n_spl_,
    g1398_p_spl_
  );


  and

  (
    g1518_p,
    g1399_n_spl_,
    g1517_n
  );


  or

  (
    g1518_n,
    g1399_p,
    g1517_p
  );


  or

  (
    g1519_n,
    g1516_p,
    g1518_n
  );


  and

  (
    g1520_p,
    n2758_lo_p_spl_001,
    lo050_buf_o2_p_spl_1
  );


  or

  (
    g1520_n,
    n2758_lo_n_spl_001,
    lo050_buf_o2_n_spl_
  );


  and

  (
    g1521_p,
    g1310_p_spl_,
    g1327_n_spl_
  );


  or

  (
    g1521_n,
    g1310_n_spl_,
    g1327_p_spl_
  );


  and

  (
    g1522_p,
    g1328_n_spl_,
    g1521_n
  );


  or

  (
    g1522_n,
    g1328_p,
    g1521_p
  );


  or

  (
    g1523_n,
    g1520_p,
    g1522_n
  );


  and

  (
    g1524_p,
    g1322_n_spl_,
    g1325_n_spl_
  );


  or

  (
    g1524_n,
    g1322_p_spl_,
    g1325_p_spl_
  );


  and

  (
    g1525_p,
    n2746_lo_p_spl_011,
    lo058_buf_o2_p_spl_1
  );


  or

  (
    g1525_n,
    n2746_lo_n_spl_011,
    lo058_buf_o2_n_spl_
  );


  and

  (
    g1526_p,
    n2734_lo_p_spl_100,
    lo062_buf_o2_p_spl_0
  );


  or

  (
    g1526_n,
    n2734_lo_n_spl_100,
    lo062_buf_o2_n_spl_0
  );


  and

  (
    g1527_p,
    g1316_n_spl_,
    g1319_n_spl_
  );


  or

  (
    g1527_n,
    g1316_p_spl_,
    g1319_p_spl_
  );


  and

  (
    g1528_p,
    g1526_n_spl_,
    g1527_n_spl_
  );


  or

  (
    g1528_n,
    g1526_p_spl_,
    g1527_p_spl_
  );


  and

  (
    g1529_p,
    g1526_p_spl_,
    g1527_p_spl_
  );


  or

  (
    g1529_n,
    g1526_n_spl_,
    g1527_n_spl_
  );


  and

  (
    g1530_p,
    g1528_n,
    g1529_n
  );


  or

  (
    g1530_n,
    g1528_p_spl_,
    g1529_p
  );


  and

  (
    g1531_p,
    g1525_n_spl_,
    g1530_p_spl_
  );


  or

  (
    g1531_n,
    g1525_p_spl_,
    g1530_n_spl_
  );


  and

  (
    g1532_p,
    g1525_p_spl_,
    g1530_n_spl_
  );


  or

  (
    g1532_n,
    g1525_n_spl_,
    g1530_p_spl_
  );


  and

  (
    g1533_p,
    g1531_n,
    g1532_n
  );


  or

  (
    g1533_n,
    g1531_p_spl_,
    g1532_p
  );


  or

  (
    g1534_n,
    g1524_p,
    g1533_n
  );


  and

  (
    g1535_p,
    g1393_n_spl_,
    g1396_n_spl_
  );


  or

  (
    g1535_n,
    g1393_p_spl_,
    g1396_p_spl_
  );


  and

  (
    g1536_p,
    n2758_lo_p_spl_010,
    lo046_buf_o2_p_spl_1
  );


  or

  (
    g1536_n,
    n2758_lo_n_spl_010,
    lo046_buf_o2_n_spl_
  );


  and

  (
    g1537_p,
    g1387_n_spl_,
    g1390_n_spl_
  );


  or

  (
    g1537_n,
    g1387_p_spl_,
    g1390_p_spl_
  );


  and

  (
    g1538_p,
    g1306_p_spl_,
    g1308_n_spl_
  );


  or

  (
    g1538_n,
    g1306_n_spl_,
    g1308_p_spl_
  );


  and

  (
    g1539_p,
    g1309_n_spl_,
    g1538_n
  );


  or

  (
    g1539_n,
    g1309_p_spl_,
    g1538_p
  );


  and

  (
    g1540_p,
    g1537_n_spl_,
    g1539_p_spl_
  );


  or

  (
    g1540_n,
    g1537_p_spl_,
    g1539_n_spl_
  );


  and

  (
    g1541_p,
    g1537_p_spl_,
    g1539_n_spl_
  );


  or

  (
    g1541_n,
    g1537_n_spl_,
    g1539_p_spl_
  );


  and

  (
    g1542_p,
    g1540_n,
    g1541_n
  );


  or

  (
    g1542_n,
    g1540_p_spl_,
    g1541_p
  );


  and

  (
    g1543_p,
    g1536_n_spl_,
    g1542_p_spl_
  );


  or

  (
    g1543_n,
    g1536_p_spl_,
    g1542_n_spl_
  );


  and

  (
    g1544_p,
    g1536_p_spl_,
    g1542_n_spl_
  );


  or

  (
    g1544_n,
    g1536_n_spl_,
    g1542_p_spl_
  );


  and

  (
    g1545_p,
    g1543_n,
    g1544_n
  );


  or

  (
    g1545_n,
    g1543_p_spl_,
    g1544_p
  );


  or

  (
    g1546_n,
    g1535_p,
    g1545_n
  );


  and

  (
    g1547_p,
    g1010_n_spl_,
    g1242_n
  );


  or

  (
    g1547_n,
    g1010_p_spl_,
    g1242_p_spl_
  );


  and

  (
    g1548_p,
    n2758_lo_p_spl_010,
    lo006_buf_o2_p_spl_0
  );


  or

  (
    g1548_n,
    n2758_lo_n_spl_010,
    lo006_buf_o2_n_spl_1
  );


  and

  (
    g1549_p,
    g1004_n_spl_,
    g1007_n_spl_
  );


  or

  (
    g1549_n,
    g1004_p_spl_,
    g1007_p_spl_
  );


  and

  (
    g1550_p,
    n2746_lo_p_spl_100,
    lo010_buf_o2_p_spl_00
  );


  or

  (
    g1550_n,
    n2746_lo_n_spl_100,
    lo010_buf_o2_n_spl_0
  );


  and

  (
    g1551_p,
    g998_n_spl_,
    g1001_n_spl_
  );


  or

  (
    g1551_n,
    g998_p_spl_,
    g1001_p_spl_
  );


  and

  (
    g1552_p,
    n2734_lo_p_spl_101,
    lo014_buf_o2_p_spl_00
  );


  or

  (
    g1552_n,
    n2734_lo_n_spl_101,
    lo014_buf_o2_n_spl_0
  );


  and

  (
    g1553_p,
    n623_o2_p,
    g995_n_spl_
  );


  or

  (
    g1553_n,
    n623_o2_n,
    g995_p_spl_
  );


  and

  (
    g1554_p,
    n655_o2_n_spl_,
    n679_o2_p_spl_
  );


  or

  (
    g1554_n,
    n655_o2_p_spl_,
    n679_o2_n_spl_
  );


  and

  (
    g1555_p,
    n655_o2_p_spl_,
    n679_o2_n_spl_
  );


  or

  (
    g1555_n,
    n655_o2_n_spl_,
    n679_o2_p_spl_
  );


  and

  (
    g1556_p,
    g1554_n_spl_,
    g1555_n
  );


  or

  (
    g1556_n,
    g1554_p_spl_,
    g1555_p
  );


  and

  (
    g1557_p,
    g1553_n_spl_,
    g1556_p_spl_
  );


  or

  (
    g1557_n,
    g1553_p_spl_,
    g1556_n_spl_
  );


  and

  (
    g1558_p,
    g1553_p_spl_,
    g1556_n_spl_
  );


  or

  (
    g1558_n,
    g1553_n_spl_,
    g1556_p_spl_
  );


  and

  (
    g1559_p,
    g1557_n_spl_,
    g1558_n
  );


  or

  (
    g1559_n,
    g1557_p_spl_,
    g1558_p
  );


  and

  (
    g1560_p,
    g1552_n_spl_,
    g1559_p_spl_
  );


  or

  (
    g1560_n,
    g1552_p_spl_,
    g1559_n_spl_
  );


  and

  (
    g1561_p,
    g1552_p_spl_,
    g1559_n_spl_
  );


  or

  (
    g1561_n,
    g1552_n_spl_,
    g1559_p_spl_
  );


  and

  (
    g1562_p,
    g1560_n_spl_,
    g1561_n
  );


  or

  (
    g1562_n,
    g1560_p_spl_,
    g1561_p
  );


  and

  (
    g1563_p,
    g1551_n_spl_,
    g1562_p_spl_
  );


  or

  (
    g1563_n,
    g1551_p_spl_,
    g1562_n_spl_
  );


  and

  (
    g1564_p,
    g1551_p_spl_,
    g1562_n_spl_
  );


  or

  (
    g1564_n,
    g1551_n_spl_,
    g1562_p_spl_
  );


  and

  (
    g1565_p,
    g1563_n_spl_,
    g1564_n
  );


  or

  (
    g1565_n,
    g1563_p_spl_,
    g1564_p
  );


  and

  (
    g1566_p,
    g1550_n_spl_,
    g1565_p_spl_
  );


  or

  (
    g1566_n,
    g1550_p_spl_,
    g1565_n_spl_
  );


  and

  (
    g1567_p,
    g1550_p_spl_,
    g1565_n_spl_
  );


  or

  (
    g1567_n,
    g1550_n_spl_,
    g1565_p_spl_
  );


  and

  (
    g1568_p,
    g1566_n_spl_,
    g1567_n
  );


  or

  (
    g1568_n,
    g1566_p_spl_,
    g1567_p
  );


  and

  (
    g1569_p,
    g1549_n_spl_,
    g1568_p_spl_
  );


  or

  (
    g1569_n,
    g1549_p_spl_,
    g1568_n_spl_
  );


  and

  (
    g1570_p,
    g1549_p_spl_,
    g1568_n_spl_
  );


  or

  (
    g1570_n,
    g1549_n_spl_,
    g1568_p_spl_
  );


  and

  (
    g1571_p,
    g1569_n_spl_,
    g1570_n
  );


  or

  (
    g1571_n,
    g1569_p_spl_,
    g1570_p
  );


  and

  (
    g1572_p,
    g1548_n_spl_,
    g1571_p_spl_
  );


  or

  (
    g1572_n,
    g1548_p_spl_,
    g1571_n_spl_
  );


  and

  (
    g1573_p,
    g1548_p_spl_,
    g1571_n_spl_
  );


  or

  (
    g1573_n,
    g1548_n_spl_,
    g1571_p_spl_
  );


  and

  (
    g1574_p,
    g1572_n_spl_,
    g1573_n
  );


  or

  (
    g1574_n,
    g1572_p_spl_,
    g1573_p
  );


  and

  (
    g1575_p,
    g1547_n_spl_,
    g1574_p_spl_
  );


  or

  (
    g1575_n,
    g1547_p,
    g1574_n
  );


  or

  (
    g1576_n,
    g1547_n_spl_,
    g1574_p_spl_
  );


  and

  (
    g1577_p,
    g1575_n,
    g1576_n
  );


  and

  (
    g1578_p,
    g1248_n_spl_,
    g1400_n
  );


  or

  (
    g1578_n,
    g1248_p_spl_,
    g1400_p_spl_
  );


  and

  (
    g1579_p,
    G2_p_spl_01,
    G19_p_spl_000
  );


  or

  (
    g1579_n,
    G2_n_spl_1,
    G19_n_spl_000
  );


  and

  (
    g1580_p,
    G4_p_spl_00,
    G17_p_spl_001
  );


  or

  (
    g1580_n,
    G4_n_spl_0,
    G17_n_spl_001
  );


  and

  (
    g1581_p,
    G3_p_spl_00,
    G18_p_spl_001
  );


  or

  (
    g1581_n,
    G3_n_spl_0,
    G18_n_spl_001
  );


  and

  (
    g1582_p,
    g1580_p_spl_,
    g1581_p_spl_
  );


  or

  (
    g1582_n,
    g1580_n_spl_,
    g1581_n_spl_
  );


  and

  (
    g1583_p,
    g1580_n_spl_,
    g1581_n_spl_
  );


  or

  (
    g1583_n,
    g1580_p_spl_,
    g1581_p_spl_
  );


  and

  (
    g1584_p,
    g1582_n_spl_0,
    g1583_n
  );


  or

  (
    g1584_n,
    g1582_p_spl_0,
    g1583_p
  );


  and

  (
    g1585_p,
    g1245_n_spl_0,
    g1584_n_spl_
  );


  or

  (
    g1585_n,
    g1245_p_spl_0,
    g1584_p_spl_
  );


  and

  (
    g1586_p,
    g1245_p_spl_,
    g1584_p_spl_
  );


  or

  (
    g1586_n,
    g1245_n_spl_,
    g1584_n_spl_
  );


  and

  (
    g1587_p,
    g1585_n_spl_,
    g1586_n
  );


  or

  (
    g1587_n,
    g1585_p_spl_,
    g1586_p
  );


  and

  (
    g1588_p,
    g1579_n_spl_,
    g1587_p_spl_
  );


  or

  (
    g1588_n,
    g1579_p_spl_,
    g1587_n_spl_
  );


  and

  (
    g1589_p,
    g1579_p_spl_,
    g1587_n_spl_
  );


  or

  (
    g1589_n,
    g1579_n_spl_,
    g1587_p_spl_
  );


  and

  (
    g1590_p,
    g1588_n_spl_,
    g1589_n
  );


  or

  (
    g1590_n,
    g1588_p_spl_,
    g1589_p
  );


  and

  (
    g1591_p,
    g1578_n_spl_,
    g1590_p_spl_
  );


  or

  (
    g1591_n,
    g1578_p,
    g1590_n
  );


  or

  (
    g1592_n,
    g1578_n_spl_,
    g1590_p_spl_
  );


  and

  (
    g1593_p,
    g1591_n,
    g1592_n
  );


  and

  (
    g1594_p,
    n2833_lo_p_spl_00,
    n6027_o2_p_spl_1
  );


  and

  (
    g1595_p,
    n2821_lo_p_spl_10,
    n6030_o2_p_spl_1
  );


  and

  (
    g1596_p,
    n2809_lo_p_spl_11,
    n6033_o2_p_spl_1
  );


  and

  (
    g1597_p,
    n2797_lo_p_spl_111,
    n6036_o2_p_spl_1
  );


  and

  (
    g1598_p,
    g1483_n_spl_,
    g1486_n_spl_
  );


  and

  (
    g1599_p,
    g1495_n_spl_,
    g1498_n_spl_
  );


  and

  (
    g1600_p,
    g1507_n_spl_,
    g1510_n_spl_
  );


  and

  (
    g1601_p,
    g1468_n_spl_,
    g1471_n_spl_
  );


  or

  (
    g1601_n,
    g1468_p_spl_,
    g1471_p_spl_
  );


  and

  (
    g1602_p,
    n2821_lo_p_spl_11,
    n6025_o2_p_spl_01
  );


  or

  (
    g1602_n,
    n2821_lo_n_spl_11,
    n6025_o2_n_spl_1
  );


  and

  (
    g1603_p,
    g1462_n_spl_,
    g1465_n_spl_
  );


  or

  (
    g1603_n,
    g1462_p_spl_,
    g1465_p_spl_
  );


  and

  (
    g1604_p,
    g1194_p_spl_,
    g1196_n_spl_
  );


  or

  (
    g1604_n,
    g1194_n_spl_,
    g1196_p_spl_
  );


  and

  (
    g1605_p,
    g1197_n_spl_,
    g1604_n
  );


  or

  (
    g1605_n,
    g1197_p_spl_,
    g1604_p
  );


  and

  (
    g1606_p,
    g1603_n_spl_,
    g1605_p_spl_
  );


  or

  (
    g1606_n,
    g1603_p_spl_,
    g1605_n_spl_
  );


  and

  (
    g1607_p,
    g1603_p_spl_,
    g1605_n_spl_
  );


  or

  (
    g1607_n,
    g1603_n_spl_,
    g1605_p_spl_
  );


  and

  (
    g1608_p,
    g1606_n_spl_,
    g1607_n
  );


  or

  (
    g1608_n,
    g1606_p_spl_,
    g1607_p
  );


  and

  (
    g1609_p,
    g1602_n_spl_,
    g1608_p_spl_
  );


  or

  (
    g1609_n,
    g1602_p_spl_,
    g1608_n_spl_
  );


  and

  (
    g1610_p,
    g1602_p_spl_,
    g1608_n_spl_
  );


  or

  (
    g1610_n,
    g1602_n_spl_,
    g1608_p_spl_
  );


  and

  (
    g1611_p,
    g1609_n_spl_,
    g1610_n
  );


  or

  (
    g1611_n,
    g1609_p_spl_,
    g1610_p
  );


  and

  (
    g1612_p,
    g1601_n_spl_,
    g1611_p_spl_
  );


  or

  (
    g1612_n,
    g1601_p_spl_,
    g1611_n_spl_
  );


  and

  (
    g1613_p,
    n2833_lo_p_spl_0,
    n6024_o2_p_spl_1
  );


  or

  (
    g1613_n,
    n2833_lo_n_spl_1,
    n6024_o2_n_spl_1
  );


  and

  (
    g1614_p,
    g1601_p_spl_,
    g1611_n_spl_
  );


  or

  (
    g1614_n,
    g1601_n_spl_,
    g1611_p_spl_
  );


  and

  (
    g1615_p,
    g1612_n_spl_,
    g1614_n
  );


  or

  (
    g1615_n,
    g1612_p,
    g1614_p
  );


  or

  (
    g1616_n,
    g1613_p,
    g1615_n
  );


  and

  (
    g1617_p,
    g1612_n_spl_,
    g1616_n_spl_
  );


  and

  (
    g1618_p,
    g1606_n_spl_,
    g1609_n_spl_
  );


  or

  (
    g1618_n,
    g1606_p_spl_,
    g1609_p_spl_
  );


  and

  (
    g1619_p,
    g1218_p_spl_,
    g1220_n_spl_
  );


  or

  (
    g1619_n,
    g1218_n_spl_,
    g1220_p_spl_
  );


  and

  (
    g1620_p,
    g1221_n_spl_,
    g1619_n
  );


  or

  (
    g1620_n,
    g1221_p_spl_,
    g1619_p
  );


  and

  (
    g1621_p,
    g1618_n_spl_,
    g1620_p_spl_
  );


  or

  (
    g1621_n,
    g1618_p_spl_,
    g1620_n_spl_
  );


  and

  (
    g1622_p,
    n2833_lo_p_spl_1,
    n6025_o2_p_spl_1
  );


  or

  (
    g1622_n,
    n2833_lo_n_spl_1,
    n6025_o2_n_spl_1
  );


  and

  (
    g1623_p,
    g1618_p_spl_,
    g1620_n_spl_
  );


  or

  (
    g1623_n,
    g1618_n_spl_,
    g1620_p_spl_
  );


  and

  (
    g1624_p,
    g1621_n_spl_,
    g1623_n
  );


  or

  (
    g1624_n,
    g1621_p,
    g1623_p
  );


  or

  (
    g1625_n,
    g1622_p,
    g1624_n
  );


  and

  (
    g1626_p,
    g1621_n_spl_,
    g1625_n_spl_
  );


  or

  (
    g1627_n,
    g1474_p,
    g1477_p_spl_
  );


  or

  (
    g1628_n,
    g1454_n_spl_,
    g1476_p_spl_
  );


  and

  (
    g1629_p,
    g1401_n_spl_,
    g1515_p_spl_
  );


  and

  (
    g1630_p,
    g1402_n_spl_,
    g1577_p_spl_
  );


  and

  (
    g1631_p,
    g1403_n_spl_,
    g1593_p_spl_
  );


  or

  (
    g1632_n,
    g1613_n,
    g1615_p
  );


  and

  (
    g1633_p,
    g1616_n_spl_,
    g1632_n
  );


  or

  (
    g1634_n,
    g1622_n,
    g1624_p
  );


  and

  (
    g1635_p,
    g1625_n_spl_,
    g1634_n
  );


  or

  (
    g1636_n,
    g1435_n,
    g1437_p
  );


  and

  (
    g1637_p,
    g1438_n_spl_,
    g1636_n
  );


  or

  (
    g1638_n,
    g1439_n,
    g1441_p
  );


  and

  (
    g1639_p,
    g1442_n_spl_,
    g1638_n
  );


  or

  (
    g1640_n,
    g1443_n,
    g1445_p
  );


  and

  (
    g1641_p,
    g1446_n_spl_,
    g1640_n
  );


  or

  (
    g1642_n,
    g1447_n,
    g1449_p
  );


  and

  (
    g1643_p,
    g1450_n_spl_,
    g1642_n
  );


  or

  (
    g1644_n,
    g1451_n,
    g1452_n
  );


  and

  (
    g1645_p,
    g1453_n_spl_,
    g1644_n
  );


  or

  (
    g1646_n,
    g1478_n,
    g1488_p
  );


  and

  (
    g1647_p,
    g1489_n_spl_,
    g1646_n
  );


  or

  (
    g1648_n,
    g1490_n,
    g1500_p
  );


  and

  (
    g1649_p,
    g1501_n_spl_,
    g1648_n
  );


  or

  (
    g1650_n,
    g1502_n,
    g1512_p
  );


  and

  (
    g1651_p,
    g1513_n_spl_,
    g1650_n
  );


  or

  (
    g1652_n,
    g1575_p,
    g1630_p_spl_
  );


  and

  (
    g1653_p,
    n2770_lo_p_spl_000,
    lo006_buf_o2_p_spl_1
  );


  or

  (
    g1653_n,
    n2770_lo_n_spl_001,
    lo006_buf_o2_n_spl_1
  );


  and

  (
    g1654_p,
    g1569_n_spl_,
    g1572_n_spl_
  );


  or

  (
    g1654_n,
    g1569_p_spl_,
    g1572_p_spl_
  );


  and

  (
    g1655_p,
    n2758_lo_p_spl_011,
    lo010_buf_o2_p_spl_0
  );


  or

  (
    g1655_n,
    n2758_lo_n_spl_011,
    lo010_buf_o2_n_spl_1
  );


  and

  (
    g1656_p,
    g1563_n_spl_,
    g1566_n_spl_
  );


  or

  (
    g1656_n,
    g1563_p_spl_,
    g1566_p_spl_
  );


  and

  (
    g1657_p,
    n2746_lo_p_spl_100,
    lo014_buf_o2_p_spl_00
  );


  or

  (
    g1657_n,
    n2746_lo_n_spl_100,
    lo014_buf_o2_n_spl_0
  );


  and

  (
    g1658_p,
    g1557_n_spl_,
    g1560_n_spl_
  );


  or

  (
    g1658_n,
    g1557_p_spl_,
    g1560_p_spl_
  );


  and

  (
    g1659_p,
    n2734_lo_p_spl_101,
    lo018_buf_o2_p_spl_00
  );


  or

  (
    g1659_n,
    n2734_lo_n_spl_101,
    lo018_buf_o2_n_spl_0
  );


  and

  (
    g1660_p,
    n677_o2_p,
    g1554_n_spl_
  );


  or

  (
    g1660_n,
    n677_o2_n,
    g1554_p_spl_
  );


  and

  (
    g1661_p,
    n717_o2_n_spl_,
    n741_o2_p_spl_
  );


  or

  (
    g1661_n,
    n717_o2_p_spl_,
    n741_o2_n_spl_
  );


  and

  (
    g1662_p,
    n717_o2_p_spl_,
    n741_o2_n_spl_
  );


  or

  (
    g1662_n,
    n717_o2_n_spl_,
    n741_o2_p_spl_
  );


  and

  (
    g1663_p,
    g1661_n_spl_,
    g1662_n
  );


  or

  (
    g1663_n,
    g1661_p_spl_,
    g1662_p
  );


  and

  (
    g1664_p,
    g1660_n_spl_,
    g1663_p_spl_
  );


  or

  (
    g1664_n,
    g1660_p_spl_,
    g1663_n_spl_
  );


  and

  (
    g1665_p,
    g1660_p_spl_,
    g1663_n_spl_
  );


  or

  (
    g1665_n,
    g1660_n_spl_,
    g1663_p_spl_
  );


  and

  (
    g1666_p,
    g1664_n_spl_,
    g1665_n
  );


  or

  (
    g1666_n,
    g1664_p_spl_,
    g1665_p
  );


  and

  (
    g1667_p,
    g1659_n_spl_,
    g1666_p_spl_
  );


  or

  (
    g1667_n,
    g1659_p_spl_,
    g1666_n_spl_
  );


  and

  (
    g1668_p,
    g1659_p_spl_,
    g1666_n_spl_
  );


  or

  (
    g1668_n,
    g1659_n_spl_,
    g1666_p_spl_
  );


  and

  (
    g1669_p,
    g1667_n_spl_,
    g1668_n
  );


  or

  (
    g1669_n,
    g1667_p_spl_,
    g1668_p
  );


  and

  (
    g1670_p,
    g1658_n_spl_,
    g1669_p_spl_
  );


  or

  (
    g1670_n,
    g1658_p_spl_,
    g1669_n_spl_
  );


  and

  (
    g1671_p,
    g1658_p_spl_,
    g1669_n_spl_
  );


  or

  (
    g1671_n,
    g1658_n_spl_,
    g1669_p_spl_
  );


  and

  (
    g1672_p,
    g1670_n_spl_,
    g1671_n
  );


  or

  (
    g1672_n,
    g1670_p_spl_,
    g1671_p
  );


  and

  (
    g1673_p,
    g1657_n_spl_,
    g1672_p_spl_
  );


  or

  (
    g1673_n,
    g1657_p_spl_,
    g1672_n_spl_
  );


  and

  (
    g1674_p,
    g1657_p_spl_,
    g1672_n_spl_
  );


  or

  (
    g1674_n,
    g1657_n_spl_,
    g1672_p_spl_
  );


  and

  (
    g1675_p,
    g1673_n_spl_,
    g1674_n
  );


  or

  (
    g1675_n,
    g1673_p_spl_,
    g1674_p
  );


  and

  (
    g1676_p,
    g1656_n_spl_,
    g1675_p_spl_
  );


  or

  (
    g1676_n,
    g1656_p_spl_,
    g1675_n_spl_
  );


  and

  (
    g1677_p,
    g1656_p_spl_,
    g1675_n_spl_
  );


  or

  (
    g1677_n,
    g1656_n_spl_,
    g1675_p_spl_
  );


  and

  (
    g1678_p,
    g1676_n_spl_,
    g1677_n
  );


  or

  (
    g1678_n,
    g1676_p_spl_,
    g1677_p
  );


  and

  (
    g1679_p,
    g1655_n_spl_,
    g1678_p_spl_
  );


  or

  (
    g1679_n,
    g1655_p_spl_,
    g1678_n_spl_
  );


  and

  (
    g1680_p,
    g1655_p_spl_,
    g1678_n_spl_
  );


  or

  (
    g1680_n,
    g1655_n_spl_,
    g1678_p_spl_
  );


  and

  (
    g1681_p,
    g1679_n_spl_,
    g1680_n
  );


  or

  (
    g1681_n,
    g1679_p_spl_,
    g1680_p
  );


  and

  (
    g1682_p,
    g1654_n_spl_,
    g1681_p_spl_
  );


  or

  (
    g1682_n,
    g1654_p_spl_,
    g1681_n_spl_
  );


  and

  (
    g1683_p,
    g1654_p_spl_,
    g1681_n_spl_
  );


  or

  (
    g1683_n,
    g1654_n_spl_,
    g1681_p_spl_
  );


  and

  (
    g1684_p,
    g1682_n_spl_,
    g1683_n
  );


  or

  (
    g1684_n,
    g1682_p,
    g1683_p
  );


  or

  (
    g1685_n,
    g1653_p,
    g1684_n
  );


  or

  (
    g1686_n,
    g1653_n,
    g1684_p
  );


  and

  (
    g1687_p,
    g1685_n_spl_,
    g1686_n
  );


  or

  (
    g1688_n,
    n2770_lo_n_spl_001,
    lo042_buf_o2_n_spl_1
  );


  or

  (
    g1689_n,
    g1535_n,
    g1545_p
  );


  and

  (
    g1690_p,
    g1546_n_spl_,
    g1689_n
  );


  and

  (
    g1691_p,
    g1688_n_spl_,
    g1690_p_spl_
  );


  or

  (
    g1692_n,
    g1688_n_spl_,
    g1690_p_spl_
  );


  or

  (
    g1693_n,
    n2758_lo_n_spl_011,
    lo054_buf_o2_n_spl_
  );


  or

  (
    g1694_n,
    g1524_n,
    g1533_p
  );


  and

  (
    g1695_p,
    g1534_n_spl_,
    g1694_n
  );


  and

  (
    g1696_p,
    g1693_n_spl_,
    g1695_p_spl_
  );


  or

  (
    g1697_n,
    g1693_n_spl_,
    g1695_p_spl_
  );


  or

  (
    g1698_n,
    n2746_lo_n_spl_101,
    lo062_buf_o2_n_spl_
  );


  or

  (
    g1699_n,
    g1528_p_spl_,
    g1531_p_spl_
  );


  and

  (
    g1700_p,
    g1698_n_spl_,
    g1699_n_spl_
  );


  or

  (
    g1701_n,
    g1698_n_spl_,
    g1699_n_spl_
  );


  or

  (
    g1702_n,
    g1540_p_spl_,
    g1543_p_spl_
  );


  or

  (
    g1703_n,
    g1520_n,
    g1522_p
  );


  and

  (
    g1704_p,
    g1523_n_spl_,
    g1703_n
  );


  and

  (
    g1705_p,
    g1702_n_spl_,
    g1704_p_spl_
  );


  or

  (
    g1706_n,
    g1702_n_spl_,
    g1704_p_spl_
  );


  and

  (
    g1707_p,
    g1676_n_spl_,
    g1679_n_spl_
  );


  or

  (
    g1707_n,
    g1676_p_spl_,
    g1679_p_spl_
  );


  and

  (
    g1708_p,
    n2758_lo_p_spl_011,
    lo014_buf_o2_p_spl_0
  );


  or

  (
    g1708_n,
    n2758_lo_n_spl_100,
    lo014_buf_o2_n_spl_1
  );


  and

  (
    g1709_p,
    g1670_n_spl_,
    g1673_n_spl_
  );


  or

  (
    g1709_n,
    g1670_p_spl_,
    g1673_p_spl_
  );


  and

  (
    g1710_p,
    n2746_lo_p_spl_101,
    lo018_buf_o2_p_spl_00
  );


  or

  (
    g1710_n,
    n2746_lo_n_spl_101,
    lo018_buf_o2_n_spl_0
  );


  and

  (
    g1711_p,
    g1664_n_spl_,
    g1667_n_spl_
  );


  or

  (
    g1711_n,
    g1664_p_spl_,
    g1667_p_spl_
  );


  and

  (
    g1712_p,
    n2734_lo_p_spl_110,
    lo022_buf_o2_p_spl_00
  );


  or

  (
    g1712_n,
    n2734_lo_n_spl_110,
    lo022_buf_o2_n_spl_0
  );


  and

  (
    g1713_p,
    n739_o2_p,
    g1661_n_spl_
  );


  or

  (
    g1713_n,
    n739_o2_n,
    g1661_p_spl_
  );


  and

  (
    g1714_p,
    n787_o2_n_spl_,
    n811_o2_p_spl_
  );


  or

  (
    g1714_n,
    n787_o2_p_spl_,
    n811_o2_n_spl_
  );


  and

  (
    g1715_p,
    n787_o2_p_spl_,
    n811_o2_n_spl_
  );


  or

  (
    g1715_n,
    n787_o2_n_spl_,
    n811_o2_p_spl_
  );


  and

  (
    g1716_p,
    g1714_n_spl_,
    g1715_n
  );


  or

  (
    g1716_n,
    g1714_p_spl_,
    g1715_p
  );


  and

  (
    g1717_p,
    g1713_n_spl_,
    g1716_p_spl_
  );


  or

  (
    g1717_n,
    g1713_p_spl_,
    g1716_n_spl_
  );


  and

  (
    g1718_p,
    g1713_p_spl_,
    g1716_n_spl_
  );


  or

  (
    g1718_n,
    g1713_n_spl_,
    g1716_p_spl_
  );


  and

  (
    g1719_p,
    g1717_n_spl_,
    g1718_n
  );


  or

  (
    g1719_n,
    g1717_p_spl_,
    g1718_p
  );


  and

  (
    g1720_p,
    g1712_n_spl_,
    g1719_p_spl_
  );


  or

  (
    g1720_n,
    g1712_p_spl_,
    g1719_n_spl_
  );


  and

  (
    g1721_p,
    g1712_p_spl_,
    g1719_n_spl_
  );


  or

  (
    g1721_n,
    g1712_n_spl_,
    g1719_p_spl_
  );


  and

  (
    g1722_p,
    g1720_n_spl_,
    g1721_n
  );


  or

  (
    g1722_n,
    g1720_p_spl_,
    g1721_p
  );


  and

  (
    g1723_p,
    g1711_n_spl_,
    g1722_p_spl_
  );


  or

  (
    g1723_n,
    g1711_p_spl_,
    g1722_n_spl_
  );


  and

  (
    g1724_p,
    g1711_p_spl_,
    g1722_n_spl_
  );


  or

  (
    g1724_n,
    g1711_n_spl_,
    g1722_p_spl_
  );


  and

  (
    g1725_p,
    g1723_n_spl_,
    g1724_n
  );


  or

  (
    g1725_n,
    g1723_p_spl_,
    g1724_p
  );


  and

  (
    g1726_p,
    g1710_n_spl_,
    g1725_p_spl_
  );


  or

  (
    g1726_n,
    g1710_p_spl_,
    g1725_n_spl_
  );


  and

  (
    g1727_p,
    g1710_p_spl_,
    g1725_n_spl_
  );


  or

  (
    g1727_n,
    g1710_n_spl_,
    g1725_p_spl_
  );


  and

  (
    g1728_p,
    g1726_n_spl_,
    g1727_n
  );


  or

  (
    g1728_n,
    g1726_p_spl_,
    g1727_p
  );


  and

  (
    g1729_p,
    g1709_n_spl_,
    g1728_p_spl_
  );


  or

  (
    g1729_n,
    g1709_p_spl_,
    g1728_n_spl_
  );


  and

  (
    g1730_p,
    g1709_p_spl_,
    g1728_n_spl_
  );


  or

  (
    g1730_n,
    g1709_n_spl_,
    g1728_p_spl_
  );


  and

  (
    g1731_p,
    g1729_n_spl_,
    g1730_n
  );


  or

  (
    g1731_n,
    g1729_p_spl_,
    g1730_p
  );


  and

  (
    g1732_p,
    g1708_n_spl_,
    g1731_p_spl_
  );


  or

  (
    g1732_n,
    g1708_p_spl_,
    g1731_n_spl_
  );


  and

  (
    g1733_p,
    g1708_p_spl_,
    g1731_n_spl_
  );


  or

  (
    g1733_n,
    g1708_n_spl_,
    g1731_p_spl_
  );


  and

  (
    g1734_p,
    g1732_n_spl_,
    g1733_n
  );


  or

  (
    g1734_n,
    g1732_p_spl_,
    g1733_p
  );


  and

  (
    g1735_p,
    g1707_n_spl_,
    g1734_p_spl_
  );


  or

  (
    g1735_n,
    g1707_p_spl_,
    g1734_n_spl_
  );


  and

  (
    g1736_p,
    n2770_lo_p_spl_001,
    lo010_buf_o2_p_spl_1
  );


  or

  (
    g1736_n,
    n2770_lo_n_spl_010,
    lo010_buf_o2_n_spl_1
  );


  and

  (
    g1737_p,
    g1707_p_spl_,
    g1734_n_spl_
  );


  or

  (
    g1737_n,
    g1707_n_spl_,
    g1734_p_spl_
  );


  and

  (
    g1738_p,
    g1735_n,
    g1737_n
  );


  or

  (
    g1738_n,
    g1735_p_spl_,
    g1737_p
  );


  and

  (
    g1739_p,
    g1736_n,
    g1738_p
  );


  or

  (
    g1740_n,
    g1735_p_spl_,
    g1739_p_spl_
  );


  and

  (
    g1741_p,
    n2770_lo_p_spl_001,
    lo014_buf_o2_p_spl_1
  );


  or

  (
    g1741_n,
    n2770_lo_n_spl_010,
    lo014_buf_o2_n_spl_1
  );


  and

  (
    g1742_p,
    g1729_n_spl_,
    g1732_n_spl_
  );


  or

  (
    g1742_n,
    g1729_p_spl_,
    g1732_p_spl_
  );


  and

  (
    g1743_p,
    n2758_lo_p_spl_100,
    lo018_buf_o2_p_spl_0
  );


  or

  (
    g1743_n,
    n2758_lo_n_spl_100,
    lo018_buf_o2_n_spl_1
  );


  and

  (
    g1744_p,
    g1723_n_spl_,
    g1726_n_spl_
  );


  or

  (
    g1744_n,
    g1723_p_spl_,
    g1726_p_spl_
  );


  and

  (
    g1745_p,
    n2746_lo_p_spl_101,
    lo022_buf_o2_p_spl_00
  );


  or

  (
    g1745_n,
    n2746_lo_n_spl_110,
    lo022_buf_o2_n_spl_0
  );


  and

  (
    g1746_p,
    g1717_n_spl_,
    g1720_n_spl_
  );


  or

  (
    g1746_n,
    g1717_p_spl_,
    g1720_p_spl_
  );


  and

  (
    g1747_p,
    n2734_lo_p_spl_110,
    lo026_buf_o2_p_spl_00
  );


  or

  (
    g1747_n,
    n2734_lo_n_spl_110,
    lo026_buf_o2_n_spl_0
  );


  and

  (
    g1748_p,
    n809_o2_p,
    g1714_n_spl_
  );


  or

  (
    g1748_n,
    n809_o2_n,
    g1714_p_spl_
  );


  and

  (
    g1749_p,
    n865_o2_n_spl_,
    n889_o2_p_spl_
  );


  or

  (
    g1749_n,
    n865_o2_p_spl_,
    n889_o2_n_spl_
  );


  and

  (
    g1750_p,
    n865_o2_p_spl_,
    n889_o2_n_spl_
  );


  or

  (
    g1750_n,
    n865_o2_n_spl_,
    n889_o2_p_spl_
  );


  and

  (
    g1751_p,
    g1749_n_spl_,
    g1750_n
  );


  or

  (
    g1751_n,
    g1749_p_spl_,
    g1750_p
  );


  and

  (
    g1752_p,
    g1748_n_spl_,
    g1751_p_spl_
  );


  or

  (
    g1752_n,
    g1748_p_spl_,
    g1751_n_spl_
  );


  and

  (
    g1753_p,
    g1748_p_spl_,
    g1751_n_spl_
  );


  or

  (
    g1753_n,
    g1748_n_spl_,
    g1751_p_spl_
  );


  and

  (
    g1754_p,
    g1752_n_spl_,
    g1753_n
  );


  or

  (
    g1754_n,
    g1752_p_spl_,
    g1753_p
  );


  and

  (
    g1755_p,
    g1747_n_spl_,
    g1754_p_spl_
  );


  or

  (
    g1755_n,
    g1747_p_spl_,
    g1754_n_spl_
  );


  and

  (
    g1756_p,
    g1747_p_spl_,
    g1754_n_spl_
  );


  or

  (
    g1756_n,
    g1747_n_spl_,
    g1754_p_spl_
  );


  and

  (
    g1757_p,
    g1755_n_spl_,
    g1756_n
  );


  or

  (
    g1757_n,
    g1755_p_spl_,
    g1756_p
  );


  and

  (
    g1758_p,
    g1746_n_spl_,
    g1757_p_spl_
  );


  or

  (
    g1758_n,
    g1746_p_spl_,
    g1757_n_spl_
  );


  and

  (
    g1759_p,
    g1746_p_spl_,
    g1757_n_spl_
  );


  or

  (
    g1759_n,
    g1746_n_spl_,
    g1757_p_spl_
  );


  and

  (
    g1760_p,
    g1758_n_spl_,
    g1759_n
  );


  or

  (
    g1760_n,
    g1758_p_spl_,
    g1759_p
  );


  and

  (
    g1761_p,
    g1745_n_spl_,
    g1760_p_spl_
  );


  or

  (
    g1761_n,
    g1745_p_spl_,
    g1760_n_spl_
  );


  and

  (
    g1762_p,
    g1745_p_spl_,
    g1760_n_spl_
  );


  or

  (
    g1762_n,
    g1745_n_spl_,
    g1760_p_spl_
  );


  and

  (
    g1763_p,
    g1761_n_spl_,
    g1762_n
  );


  or

  (
    g1763_n,
    g1761_p_spl_,
    g1762_p
  );


  and

  (
    g1764_p,
    g1744_n_spl_,
    g1763_p_spl_
  );


  or

  (
    g1764_n,
    g1744_p_spl_,
    g1763_n_spl_
  );


  and

  (
    g1765_p,
    g1744_p_spl_,
    g1763_n_spl_
  );


  or

  (
    g1765_n,
    g1744_n_spl_,
    g1763_p_spl_
  );


  and

  (
    g1766_p,
    g1764_n_spl_,
    g1765_n
  );


  or

  (
    g1766_n,
    g1764_p_spl_,
    g1765_p
  );


  and

  (
    g1767_p,
    g1743_n_spl_,
    g1766_p_spl_
  );


  or

  (
    g1767_n,
    g1743_p_spl_,
    g1766_n_spl_
  );


  and

  (
    g1768_p,
    g1743_p_spl_,
    g1766_n_spl_
  );


  or

  (
    g1768_n,
    g1743_n_spl_,
    g1766_p_spl_
  );


  and

  (
    g1769_p,
    g1767_n_spl_,
    g1768_n
  );


  or

  (
    g1769_n,
    g1767_p_spl_,
    g1768_p
  );


  and

  (
    g1770_p,
    g1742_n_spl_,
    g1769_p_spl_
  );


  or

  (
    g1770_n,
    g1742_p_spl_,
    g1769_n_spl_
  );


  and

  (
    g1771_p,
    g1742_p_spl_,
    g1769_n_spl_
  );


  or

  (
    g1771_n,
    g1742_n_spl_,
    g1769_p_spl_
  );


  and

  (
    g1772_p,
    g1770_n,
    g1771_n
  );


  or

  (
    g1772_n,
    g1770_p_spl_,
    g1771_p
  );


  and

  (
    g1773_p,
    g1741_n_spl_,
    g1772_p_spl_
  );


  or

  (
    g1773_n,
    g1741_p,
    g1772_n
  );


  or

  (
    g1774_n,
    g1741_n_spl_,
    g1772_p_spl_
  );


  and

  (
    g1775_p,
    g1773_n,
    g1774_n
  );


  and

  (
    g1776_p,
    g1740_n_spl_,
    g1775_p_spl_
  );


  or

  (
    g1777_n,
    g1740_n_spl_,
    g1775_p_spl_
  );


  or

  (
    g1778_n,
    g1770_p_spl_,
    g1773_p
  );


  and

  (
    g1779_p,
    n2770_lo_p_spl_01,
    lo018_buf_o2_p_spl_1
  );


  or

  (
    g1779_n,
    n2770_lo_n_spl_01,
    lo018_buf_o2_n_spl_1
  );


  and

  (
    g1780_p,
    g1764_n_spl_,
    g1767_n_spl_
  );


  or

  (
    g1780_n,
    g1764_p_spl_,
    g1767_p_spl_
  );


  and

  (
    g1781_p,
    n2758_lo_p_spl_100,
    lo022_buf_o2_p_spl_0
  );


  or

  (
    g1781_n,
    n2758_lo_n_spl_101,
    lo022_buf_o2_n_spl_1
  );


  and

  (
    g1782_p,
    g1758_n_spl_,
    g1761_n_spl_
  );


  or

  (
    g1782_n,
    g1758_p_spl_,
    g1761_p_spl_
  );


  and

  (
    g1783_p,
    n2746_lo_p_spl_110,
    lo026_buf_o2_p_spl_00
  );


  or

  (
    g1783_n,
    n2746_lo_n_spl_110,
    lo026_buf_o2_n_spl_0
  );


  and

  (
    g1784_p,
    g1752_n_spl_,
    g1755_n_spl_
  );


  or

  (
    g1784_n,
    g1752_p_spl_,
    g1755_p_spl_
  );


  and

  (
    g1785_p,
    n2734_lo_p_spl_111,
    lo030_buf_o2_p_spl_00
  );


  or

  (
    g1785_n,
    n2734_lo_n_spl_111,
    lo030_buf_o2_n_spl_0
  );


  and

  (
    g1786_p,
    n887_o2_p,
    g1749_n_spl_
  );


  or

  (
    g1786_n,
    n887_o2_n,
    g1749_p_spl_
  );


  and

  (
    g1787_p,
    n951_o2_n_spl_,
    n975_o2_p_spl_
  );


  or

  (
    g1787_n,
    n951_o2_p_spl_,
    n975_o2_n_spl_
  );


  and

  (
    g1788_p,
    n951_o2_p_spl_,
    n975_o2_n_spl_
  );


  or

  (
    g1788_n,
    n951_o2_n_spl_,
    n975_o2_p_spl_
  );


  and

  (
    g1789_p,
    g1787_n_spl_,
    g1788_n
  );


  or

  (
    g1789_n,
    g1787_p_spl_,
    g1788_p
  );


  and

  (
    g1790_p,
    g1786_n_spl_,
    g1789_p_spl_
  );


  or

  (
    g1790_n,
    g1786_p_spl_,
    g1789_n_spl_
  );


  and

  (
    g1791_p,
    g1786_p_spl_,
    g1789_n_spl_
  );


  or

  (
    g1791_n,
    g1786_n_spl_,
    g1789_p_spl_
  );


  and

  (
    g1792_p,
    g1790_n_spl_,
    g1791_n
  );


  or

  (
    g1792_n,
    g1790_p_spl_,
    g1791_p
  );


  and

  (
    g1793_p,
    g1785_n_spl_,
    g1792_p_spl_
  );


  or

  (
    g1793_n,
    g1785_p_spl_,
    g1792_n_spl_
  );


  and

  (
    g1794_p,
    g1785_p_spl_,
    g1792_n_spl_
  );


  or

  (
    g1794_n,
    g1785_n_spl_,
    g1792_p_spl_
  );


  and

  (
    g1795_p,
    g1793_n_spl_,
    g1794_n
  );


  or

  (
    g1795_n,
    g1793_p_spl_,
    g1794_p
  );


  and

  (
    g1796_p,
    g1784_n_spl_,
    g1795_p_spl_
  );


  or

  (
    g1796_n,
    g1784_p_spl_,
    g1795_n_spl_
  );


  and

  (
    g1797_p,
    g1784_p_spl_,
    g1795_n_spl_
  );


  or

  (
    g1797_n,
    g1784_n_spl_,
    g1795_p_spl_
  );


  and

  (
    g1798_p,
    g1796_n_spl_,
    g1797_n
  );


  or

  (
    g1798_n,
    g1796_p_spl_,
    g1797_p
  );


  and

  (
    g1799_p,
    g1783_n_spl_,
    g1798_p_spl_
  );


  or

  (
    g1799_n,
    g1783_p_spl_,
    g1798_n_spl_
  );


  and

  (
    g1800_p,
    g1783_p_spl_,
    g1798_n_spl_
  );


  or

  (
    g1800_n,
    g1783_n_spl_,
    g1798_p_spl_
  );


  and

  (
    g1801_p,
    g1799_n_spl_,
    g1800_n
  );


  or

  (
    g1801_n,
    g1799_p_spl_,
    g1800_p
  );


  and

  (
    g1802_p,
    g1782_n_spl_,
    g1801_p_spl_
  );


  or

  (
    g1802_n,
    g1782_p_spl_,
    g1801_n_spl_
  );


  and

  (
    g1803_p,
    g1782_p_spl_,
    g1801_n_spl_
  );


  or

  (
    g1803_n,
    g1782_n_spl_,
    g1801_p_spl_
  );


  and

  (
    g1804_p,
    g1802_n_spl_,
    g1803_n
  );


  or

  (
    g1804_n,
    g1802_p_spl_,
    g1803_p
  );


  and

  (
    g1805_p,
    g1781_n_spl_,
    g1804_p_spl_
  );


  or

  (
    g1805_n,
    g1781_p_spl_,
    g1804_n_spl_
  );


  and

  (
    g1806_p,
    g1781_p_spl_,
    g1804_n_spl_
  );


  or

  (
    g1806_n,
    g1781_n_spl_,
    g1804_p_spl_
  );


  and

  (
    g1807_p,
    g1805_n_spl_,
    g1806_n
  );


  or

  (
    g1807_n,
    g1805_p_spl_,
    g1806_p
  );


  and

  (
    g1808_p,
    g1780_n_spl_,
    g1807_p_spl_
  );


  or

  (
    g1808_n,
    g1780_p_spl_,
    g1807_n_spl_
  );


  and

  (
    g1809_p,
    g1780_p_spl_,
    g1807_n_spl_
  );


  or

  (
    g1809_n,
    g1780_n_spl_,
    g1807_p_spl_
  );


  and

  (
    g1810_p,
    g1808_n,
    g1809_n
  );


  or

  (
    g1810_n,
    g1808_p_spl_,
    g1809_p
  );


  and

  (
    g1811_p,
    g1779_n_spl_,
    g1810_p_spl_
  );


  or

  (
    g1811_n,
    g1779_p,
    g1810_n
  );


  or

  (
    g1812_n,
    g1779_n_spl_,
    g1810_p_spl_
  );


  and

  (
    g1813_p,
    g1811_n,
    g1812_n
  );


  and

  (
    g1814_p,
    g1778_n_spl_,
    g1813_p_spl_
  );


  or

  (
    g1815_n,
    g1778_n_spl_,
    g1813_p_spl_
  );


  or

  (
    g1816_n,
    g1808_p_spl_,
    g1811_p
  );


  and

  (
    g1817_p,
    n2770_lo_p_spl_01,
    lo022_buf_o2_p_spl_1
  );


  or

  (
    g1817_n,
    n2770_lo_n_spl_10,
    lo022_buf_o2_n_spl_1
  );


  and

  (
    g1818_p,
    g1802_n_spl_,
    g1805_n_spl_
  );


  or

  (
    g1818_n,
    g1802_p_spl_,
    g1805_p_spl_
  );


  and

  (
    g1819_p,
    n2758_lo_p_spl_101,
    lo026_buf_o2_p_spl_0
  );


  or

  (
    g1819_n,
    n2758_lo_n_spl_101,
    lo026_buf_o2_n_spl_1
  );


  and

  (
    g1820_p,
    g1796_n_spl_,
    g1799_n_spl_
  );


  or

  (
    g1820_n,
    g1796_p_spl_,
    g1799_p_spl_
  );


  and

  (
    g1821_p,
    n2746_lo_p_spl_110,
    lo030_buf_o2_p_spl_00
  );


  or

  (
    g1821_n,
    n2746_lo_n_spl_111,
    lo030_buf_o2_n_spl_0
  );


  and

  (
    g1822_p,
    g1790_n_spl_,
    g1793_n_spl_
  );


  or

  (
    g1822_n,
    g1790_p_spl_,
    g1793_p_spl_
  );


  and

  (
    g1823_p,
    n2734_lo_p_spl_111,
    lo034_buf_o2_p_spl_00
  );


  or

  (
    g1823_n,
    n2734_lo_n_spl_111,
    lo034_buf_o2_n_spl_0
  );


  and

  (
    g1824_p,
    n973_o2_p,
    g1787_n_spl_
  );


  or

  (
    g1824_n,
    n973_o2_n,
    g1787_p_spl_
  );


  and

  (
    g1825_p,
    n1045_o2_p_spl_,
    n1069_o2_n_spl_
  );


  or

  (
    g1825_n,
    n1045_o2_n_spl_,
    n1069_o2_p_spl_
  );


  and

  (
    g1826_p,
    g1329_n_spl_,
    g1825_n
  );


  or

  (
    g1826_n,
    g1329_p_spl_,
    g1825_p
  );


  and

  (
    g1827_p,
    g1824_n_spl_,
    g1826_p_spl_
  );


  or

  (
    g1827_n,
    g1824_p_spl_,
    g1826_n_spl_
  );


  and

  (
    g1828_p,
    g1824_p_spl_,
    g1826_n_spl_
  );


  or

  (
    g1828_n,
    g1824_n_spl_,
    g1826_p_spl_
  );


  and

  (
    g1829_p,
    g1827_n_spl_,
    g1828_n
  );


  or

  (
    g1829_n,
    g1827_p_spl_,
    g1828_p
  );


  and

  (
    g1830_p,
    g1823_n_spl_,
    g1829_p_spl_
  );


  or

  (
    g1830_n,
    g1823_p_spl_,
    g1829_n_spl_
  );


  and

  (
    g1831_p,
    g1823_p_spl_,
    g1829_n_spl_
  );


  or

  (
    g1831_n,
    g1823_n_spl_,
    g1829_p_spl_
  );


  and

  (
    g1832_p,
    g1830_n_spl_,
    g1831_n
  );


  or

  (
    g1832_n,
    g1830_p_spl_,
    g1831_p
  );


  and

  (
    g1833_p,
    g1822_n_spl_,
    g1832_p_spl_
  );


  or

  (
    g1833_n,
    g1822_p_spl_,
    g1832_n_spl_
  );


  and

  (
    g1834_p,
    g1822_p_spl_,
    g1832_n_spl_
  );


  or

  (
    g1834_n,
    g1822_n_spl_,
    g1832_p_spl_
  );


  and

  (
    g1835_p,
    g1833_n_spl_,
    g1834_n
  );


  or

  (
    g1835_n,
    g1833_p_spl_,
    g1834_p
  );


  and

  (
    g1836_p,
    g1821_n_spl_,
    g1835_p_spl_
  );


  or

  (
    g1836_n,
    g1821_p_spl_,
    g1835_n_spl_
  );


  and

  (
    g1837_p,
    g1821_p_spl_,
    g1835_n_spl_
  );


  or

  (
    g1837_n,
    g1821_n_spl_,
    g1835_p_spl_
  );


  and

  (
    g1838_p,
    g1836_n_spl_,
    g1837_n
  );


  or

  (
    g1838_n,
    g1836_p_spl_,
    g1837_p
  );


  and

  (
    g1839_p,
    g1820_n_spl_,
    g1838_p_spl_
  );


  or

  (
    g1839_n,
    g1820_p_spl_,
    g1838_n_spl_
  );


  and

  (
    g1840_p,
    g1820_p_spl_,
    g1838_n_spl_
  );


  or

  (
    g1840_n,
    g1820_n_spl_,
    g1838_p_spl_
  );


  and

  (
    g1841_p,
    g1839_n_spl_,
    g1840_n
  );


  or

  (
    g1841_n,
    g1839_p_spl_,
    g1840_p
  );


  and

  (
    g1842_p,
    g1819_n_spl_,
    g1841_p_spl_
  );


  or

  (
    g1842_n,
    g1819_p_spl_,
    g1841_n_spl_
  );


  and

  (
    g1843_p,
    g1819_p_spl_,
    g1841_n_spl_
  );


  or

  (
    g1843_n,
    g1819_n_spl_,
    g1841_p_spl_
  );


  and

  (
    g1844_p,
    g1842_n_spl_,
    g1843_n
  );


  or

  (
    g1844_n,
    g1842_p_spl_,
    g1843_p
  );


  and

  (
    g1845_p,
    g1818_n_spl_,
    g1844_p_spl_
  );


  or

  (
    g1845_n,
    g1818_p_spl_,
    g1844_n_spl_
  );


  and

  (
    g1846_p,
    g1818_p_spl_,
    g1844_n_spl_
  );


  or

  (
    g1846_n,
    g1818_n_spl_,
    g1844_p_spl_
  );


  and

  (
    g1847_p,
    g1845_n,
    g1846_n
  );


  or

  (
    g1847_n,
    g1845_p_spl_,
    g1846_p
  );


  and

  (
    g1848_p,
    g1817_n_spl_,
    g1847_p_spl_
  );


  or

  (
    g1848_n,
    g1817_p,
    g1847_n
  );


  or

  (
    g1849_n,
    g1817_n_spl_,
    g1847_p_spl_
  );


  and

  (
    g1850_p,
    g1848_n,
    g1849_n
  );


  and

  (
    g1851_p,
    g1816_n_spl_,
    g1850_p_spl_
  );


  or

  (
    g1852_n,
    g1816_n_spl_,
    g1850_p_spl_
  );


  or

  (
    g1853_n,
    g1845_p_spl_,
    g1848_p
  );


  and

  (
    g1854_p,
    n2770_lo_p_spl_10,
    lo026_buf_o2_p_spl_1
  );


  or

  (
    g1854_n,
    n2770_lo_n_spl_10,
    lo026_buf_o2_n_spl_1
  );


  and

  (
    g1855_p,
    g1839_n_spl_,
    g1842_n_spl_
  );


  or

  (
    g1855_n,
    g1839_p_spl_,
    g1842_p_spl_
  );


  and

  (
    g1856_p,
    n2758_lo_p_spl_101,
    lo030_buf_o2_p_spl_0
  );


  or

  (
    g1856_n,
    n2758_lo_n_spl_11,
    lo030_buf_o2_n_spl_1
  );


  and

  (
    g1857_p,
    g1833_n_spl_,
    g1836_n_spl_
  );


  or

  (
    g1857_n,
    g1833_p_spl_,
    g1836_p_spl_
  );


  and

  (
    g1858_p,
    n2746_lo_p_spl_11,
    lo034_buf_o2_p_spl_00
  );


  or

  (
    g1858_n,
    n2746_lo_n_spl_111,
    lo034_buf_o2_n_spl_0
  );


  and

  (
    g1859_p,
    g1827_n_spl_,
    g1830_n_spl_
  );


  or

  (
    g1859_n,
    g1827_p_spl_,
    g1830_p_spl_
  );


  and

  (
    g1860_p,
    g1335_p_spl_,
    g1337_n_spl_
  );


  or

  (
    g1860_n,
    g1335_n_spl_,
    g1337_p_spl_
  );


  and

  (
    g1861_p,
    g1338_n_spl_,
    g1860_n
  );


  or

  (
    g1861_n,
    g1338_p_spl_,
    g1860_p
  );


  and

  (
    g1862_p,
    g1859_n_spl_,
    g1861_p_spl_
  );


  or

  (
    g1862_n,
    g1859_p_spl_,
    g1861_n_spl_
  );


  and

  (
    g1863_p,
    g1859_p_spl_,
    g1861_n_spl_
  );


  or

  (
    g1863_n,
    g1859_n_spl_,
    g1861_p_spl_
  );


  and

  (
    g1864_p,
    g1862_n_spl_,
    g1863_n
  );


  or

  (
    g1864_n,
    g1862_p_spl_,
    g1863_p
  );


  and

  (
    g1865_p,
    g1858_n_spl_,
    g1864_p_spl_
  );


  or

  (
    g1865_n,
    g1858_p_spl_,
    g1864_n_spl_
  );


  and

  (
    g1866_p,
    g1858_p_spl_,
    g1864_n_spl_
  );


  or

  (
    g1866_n,
    g1858_n_spl_,
    g1864_p_spl_
  );


  and

  (
    g1867_p,
    g1865_n_spl_,
    g1866_n
  );


  or

  (
    g1867_n,
    g1865_p_spl_,
    g1866_p
  );


  and

  (
    g1868_p,
    g1857_n_spl_,
    g1867_p_spl_
  );


  or

  (
    g1868_n,
    g1857_p_spl_,
    g1867_n_spl_
  );


  and

  (
    g1869_p,
    g1857_p_spl_,
    g1867_n_spl_
  );


  or

  (
    g1869_n,
    g1857_n_spl_,
    g1867_p_spl_
  );


  and

  (
    g1870_p,
    g1868_n_spl_,
    g1869_n
  );


  or

  (
    g1870_n,
    g1868_p_spl_,
    g1869_p
  );


  and

  (
    g1871_p,
    g1856_n_spl_,
    g1870_p_spl_
  );


  or

  (
    g1871_n,
    g1856_p_spl_,
    g1870_n_spl_
  );


  and

  (
    g1872_p,
    g1856_p_spl_,
    g1870_n_spl_
  );


  or

  (
    g1872_n,
    g1856_n_spl_,
    g1870_p_spl_
  );


  and

  (
    g1873_p,
    g1871_n_spl_,
    g1872_n
  );


  or

  (
    g1873_n,
    g1871_p_spl_,
    g1872_p
  );


  and

  (
    g1874_p,
    g1855_n_spl_,
    g1873_p_spl_
  );


  or

  (
    g1874_n,
    g1855_p_spl_,
    g1873_n_spl_
  );


  and

  (
    g1875_p,
    g1855_p_spl_,
    g1873_n_spl_
  );


  or

  (
    g1875_n,
    g1855_n_spl_,
    g1873_p_spl_
  );


  and

  (
    g1876_p,
    g1874_n,
    g1875_n
  );


  or

  (
    g1876_n,
    g1874_p_spl_,
    g1875_p
  );


  and

  (
    g1877_p,
    g1854_n_spl_,
    g1876_p_spl_
  );


  or

  (
    g1877_n,
    g1854_p,
    g1876_n
  );


  or

  (
    g1878_n,
    g1854_n_spl_,
    g1876_p_spl_
  );


  and

  (
    g1879_p,
    g1877_n,
    g1878_n
  );


  and

  (
    g1880_p,
    g1853_n_spl_,
    g1879_p_spl_
  );


  or

  (
    g1881_n,
    g1853_n_spl_,
    g1879_p_spl_
  );


  or

  (
    g1882_n,
    g1874_p_spl_,
    g1877_p
  );


  and

  (
    g1883_p,
    n2770_lo_p_spl_10,
    lo030_buf_o2_p_spl_1
  );


  or

  (
    g1883_n,
    n2770_lo_n_spl_11,
    lo030_buf_o2_n_spl_1
  );


  and

  (
    g1884_p,
    g1868_n_spl_,
    g1871_n_spl_
  );


  or

  (
    g1884_n,
    g1868_p_spl_,
    g1871_p_spl_
  );


  and

  (
    g1885_p,
    n2758_lo_p_spl_11,
    lo034_buf_o2_p_spl_0
  );


  or

  (
    g1885_n,
    n2758_lo_n_spl_11,
    lo034_buf_o2_n_spl_1
  );


  and

  (
    g1886_p,
    g1862_n_spl_,
    g1865_n_spl_
  );


  or

  (
    g1886_n,
    g1862_p_spl_,
    g1865_p_spl_
  );


  and

  (
    g1887_p,
    g1352_p_spl_,
    g1354_n_spl_
  );


  or

  (
    g1887_n,
    g1352_n_spl_,
    g1354_p_spl_
  );


  and

  (
    g1888_p,
    g1355_n_spl_,
    g1887_n
  );


  or

  (
    g1888_n,
    g1355_p_spl_,
    g1887_p
  );


  and

  (
    g1889_p,
    g1886_n_spl_,
    g1888_p_spl_
  );


  or

  (
    g1889_n,
    g1886_p_spl_,
    g1888_n_spl_
  );


  and

  (
    g1890_p,
    g1886_p_spl_,
    g1888_n_spl_
  );


  or

  (
    g1890_n,
    g1886_n_spl_,
    g1888_p_spl_
  );


  and

  (
    g1891_p,
    g1889_n_spl_,
    g1890_n
  );


  or

  (
    g1891_n,
    g1889_p_spl_,
    g1890_p
  );


  and

  (
    g1892_p,
    g1885_n_spl_,
    g1891_p_spl_
  );


  or

  (
    g1892_n,
    g1885_p_spl_,
    g1891_n_spl_
  );


  and

  (
    g1893_p,
    g1885_p_spl_,
    g1891_n_spl_
  );


  or

  (
    g1893_n,
    g1885_n_spl_,
    g1891_p_spl_
  );


  and

  (
    g1894_p,
    g1892_n_spl_,
    g1893_n
  );


  or

  (
    g1894_n,
    g1892_p_spl_,
    g1893_p
  );


  and

  (
    g1895_p,
    g1884_n_spl_,
    g1894_p_spl_
  );


  or

  (
    g1895_n,
    g1884_p_spl_,
    g1894_n_spl_
  );


  and

  (
    g1896_p,
    g1884_p_spl_,
    g1894_n_spl_
  );


  or

  (
    g1896_n,
    g1884_n_spl_,
    g1894_p_spl_
  );


  and

  (
    g1897_p,
    g1895_n,
    g1896_n
  );


  or

  (
    g1897_n,
    g1895_p_spl_,
    g1896_p
  );


  and

  (
    g1898_p,
    g1883_n_spl_,
    g1897_p_spl_
  );


  or

  (
    g1898_n,
    g1883_p,
    g1897_n
  );


  or

  (
    g1899_n,
    g1883_n_spl_,
    g1897_p_spl_
  );


  and

  (
    g1900_p,
    g1898_n,
    g1899_n
  );


  and

  (
    g1901_p,
    g1882_n_spl_,
    g1900_p_spl_
  );


  or

  (
    g1902_n,
    g1882_n_spl_,
    g1900_p_spl_
  );


  or

  (
    g1903_n,
    g1895_p_spl_,
    g1898_p
  );


  and

  (
    g1904_p,
    n2770_lo_p_spl_11,
    lo034_buf_o2_p_spl_1
  );


  or

  (
    g1904_n,
    n2770_lo_n_spl_11,
    lo034_buf_o2_n_spl_1
  );


  and

  (
    g1905_p,
    g1889_n_spl_,
    g1892_n_spl_
  );


  or

  (
    g1905_n,
    g1889_p_spl_,
    g1892_p_spl_
  );


  and

  (
    g1906_p,
    g1376_p_spl_,
    g1378_n_spl_
  );


  or

  (
    g1906_n,
    g1376_n_spl_,
    g1378_p_spl_
  );


  and

  (
    g1907_p,
    g1379_n_spl_,
    g1906_n
  );


  or

  (
    g1907_n,
    g1379_p_spl_,
    g1906_p
  );


  and

  (
    g1908_p,
    g1905_n_spl_,
    g1907_p_spl_
  );


  or

  (
    g1908_n,
    g1905_p_spl_,
    g1907_n_spl_
  );


  and

  (
    g1909_p,
    g1905_p_spl_,
    g1907_n_spl_
  );


  or

  (
    g1909_n,
    g1905_n_spl_,
    g1907_p_spl_
  );


  and

  (
    g1910_p,
    g1908_n,
    g1909_n
  );


  or

  (
    g1910_n,
    g1908_p_spl_,
    g1909_p
  );


  and

  (
    g1911_p,
    g1904_n_spl_,
    g1910_p_spl_
  );


  or

  (
    g1911_n,
    g1904_p,
    g1910_n
  );


  or

  (
    g1912_n,
    g1904_n_spl_,
    g1910_p_spl_
  );


  and

  (
    g1913_p,
    g1911_n,
    g1912_n
  );


  and

  (
    g1914_p,
    g1903_n_spl_,
    g1913_p_spl_
  );


  or

  (
    g1915_n,
    g1903_n_spl_,
    g1913_p_spl_
  );


  or

  (
    g1916_n,
    g1908_p_spl_,
    g1911_p
  );


  or

  (
    g1917_n,
    g1516_n,
    g1518_p
  );


  and

  (
    g1918_p,
    g1519_n_spl_,
    g1917_n
  );


  and

  (
    g1919_p,
    g1916_n_spl_,
    g1918_p_spl_
  );


  or

  (
    g1920_n,
    g1916_n_spl_,
    g1918_p_spl_
  );


  and

  (
    g1921_p,
    g1682_n_spl_,
    g1685_n_spl_
  );


  and

  (
    g1922_p,
    g1736_p,
    g1738_n
  );


  or

  (
    g1923_n,
    g1739_p_spl_,
    g1922_p
  );


  or

  (
    g1924_n,
    g1921_p_spl_,
    g1923_n_spl_
  );


  and

  (
    g1925_p,
    g1921_p_spl_,
    g1923_n_spl_
  );


  and

  (
    g1926_p,
    G5_p_spl_00,
    G17_p_spl_001
  );


  or

  (
    g1926_n,
    G5_n_spl_0,
    G17_n_spl_001
  );


  and

  (
    g1927_p,
    G4_p_spl_00,
    G18_p_spl_001
  );


  or

  (
    g1927_n,
    G4_n_spl_0,
    G18_n_spl_001
  );


  and

  (
    g1928_p,
    g1926_p_spl_,
    g1927_p_spl_
  );


  or

  (
    g1928_n,
    g1926_n_spl_,
    g1927_n_spl_
  );


  and

  (
    g1929_p,
    g1926_n_spl_,
    g1927_n_spl_
  );


  or

  (
    g1929_n,
    g1926_p_spl_,
    g1927_p_spl_
  );


  and

  (
    g1930_p,
    g1928_n_spl_0,
    g1929_n
  );


  or

  (
    g1930_n,
    g1928_p_spl_0,
    g1929_p
  );


  and

  (
    g1931_p,
    g1582_n_spl_0,
    g1930_n_spl_
  );


  or

  (
    g1931_n,
    g1582_p_spl_0,
    g1930_p_spl_
  );


  and

  (
    g1932_p,
    G3_p_spl_01,
    G19_p_spl_001
  );


  or

  (
    g1932_n,
    G3_n_spl_1,
    G19_n_spl_001
  );


  and

  (
    g1933_p,
    g1582_p_spl_,
    g1930_p_spl_
  );


  or

  (
    g1933_n,
    g1582_n_spl_,
    g1930_n_spl_
  );


  and

  (
    g1934_p,
    g1931_n_spl_,
    g1933_n
  );


  or

  (
    g1934_n,
    g1931_p_spl_,
    g1933_p
  );


  and

  (
    g1935_p,
    g1932_n_spl_,
    g1934_p_spl_
  );


  or

  (
    g1935_n,
    g1932_p_spl_,
    g1934_n_spl_
  );


  and

  (
    g1936_p,
    g1931_n_spl_,
    g1935_n_spl_
  );


  or

  (
    g1936_n,
    g1931_p_spl_,
    g1935_p_spl_
  );


  and

  (
    g1937_p,
    G4_p_spl_01,
    G19_p_spl_001
  );


  or

  (
    g1937_n,
    G4_n_spl_1,
    G19_n_spl_001
  );


  and

  (
    g1938_p,
    G6_p_spl_00,
    G17_p_spl_010
  );


  or

  (
    g1938_n,
    G6_n_spl_0,
    G17_n_spl_010
  );


  and

  (
    g1939_p,
    G5_p_spl_00,
    G18_p_spl_010
  );


  or

  (
    g1939_n,
    G5_n_spl_0,
    G18_n_spl_010
  );


  and

  (
    g1940_p,
    g1938_p_spl_,
    g1939_p_spl_
  );


  or

  (
    g1940_n,
    g1938_n_spl_,
    g1939_n_spl_
  );


  and

  (
    g1941_p,
    g1938_n_spl_,
    g1939_n_spl_
  );


  or

  (
    g1941_n,
    g1938_p_spl_,
    g1939_p_spl_
  );


  and

  (
    g1942_p,
    g1940_n_spl_0,
    g1941_n
  );


  or

  (
    g1942_n,
    g1940_p_spl_0,
    g1941_p
  );


  and

  (
    g1943_p,
    g1928_n_spl_0,
    g1942_n_spl_
  );


  or

  (
    g1943_n,
    g1928_p_spl_0,
    g1942_p_spl_
  );


  and

  (
    g1944_p,
    g1928_p_spl_,
    g1942_p_spl_
  );


  or

  (
    g1944_n,
    g1928_n_spl_,
    g1942_n_spl_
  );


  and

  (
    g1945_p,
    g1943_n_spl_,
    g1944_n
  );


  or

  (
    g1945_n,
    g1943_p_spl_,
    g1944_p
  );


  and

  (
    g1946_p,
    g1937_n_spl_,
    g1945_p_spl_
  );


  or

  (
    g1946_n,
    g1937_p_spl_,
    g1945_n_spl_
  );


  and

  (
    g1947_p,
    g1937_p_spl_,
    g1945_n_spl_
  );


  or

  (
    g1947_n,
    g1937_n_spl_,
    g1945_p_spl_
  );


  and

  (
    g1948_p,
    g1946_n_spl_,
    g1947_n
  );


  or

  (
    g1948_n,
    g1946_p_spl_,
    g1947_p
  );


  and

  (
    g1949_p,
    g1936_n_spl_,
    g1948_p_spl_
  );


  or

  (
    g1949_n,
    g1936_p_spl_,
    g1948_n_spl_
  );


  and

  (
    g1950_p,
    G3_p_spl_01,
    G20_p_spl_000
  );


  or

  (
    g1950_n,
    G3_n_spl_1,
    G20_n_spl_000
  );


  and

  (
    g1951_p,
    g1936_p_spl_,
    g1948_n_spl_
  );


  or

  (
    g1951_n,
    g1936_n_spl_,
    g1948_p_spl_
  );


  and

  (
    g1952_p,
    g1949_n_spl_,
    g1951_n
  );


  or

  (
    g1952_n,
    g1949_p_spl_,
    g1951_p
  );


  and

  (
    g1953_p,
    g1950_n_spl_,
    g1952_p_spl_
  );


  or

  (
    g1953_n,
    g1950_p_spl_,
    g1952_n_spl_
  );


  and

  (
    g1954_p,
    g1949_n_spl_,
    g1953_n_spl_
  );


  or

  (
    g1954_n,
    g1949_p_spl_,
    g1953_p_spl_
  );


  and

  (
    g1955_p,
    G4_p_spl_01,
    G20_p_spl_000
  );


  or

  (
    g1955_n,
    G4_n_spl_1,
    G20_n_spl_001
  );


  and

  (
    g1956_p,
    g1943_n_spl_,
    g1946_n_spl_
  );


  or

  (
    g1956_n,
    g1943_p_spl_,
    g1946_p_spl_
  );


  and

  (
    g1957_p,
    G5_p_spl_01,
    G19_p_spl_010
  );


  or

  (
    g1957_n,
    G5_n_spl_1,
    G19_n_spl_010
  );


  and

  (
    g1958_p,
    G7_p_spl_00,
    G17_p_spl_010
  );


  or

  (
    g1958_n,
    G7_n_spl_0,
    G17_n_spl_010
  );


  and

  (
    g1959_p,
    G6_p_spl_00,
    G18_p_spl_010
  );


  or

  (
    g1959_n,
    G6_n_spl_0,
    G18_n_spl_010
  );


  and

  (
    g1960_p,
    g1958_p_spl_,
    g1959_p_spl_
  );


  or

  (
    g1960_n,
    g1958_n_spl_,
    g1959_n_spl_
  );


  and

  (
    g1961_p,
    g1958_n_spl_,
    g1959_n_spl_
  );


  or

  (
    g1961_n,
    g1958_p_spl_,
    g1959_p_spl_
  );


  and

  (
    g1962_p,
    g1960_n_spl_0,
    g1961_n
  );


  or

  (
    g1962_n,
    g1960_p_spl_0,
    g1961_p
  );


  and

  (
    g1963_p,
    g1940_n_spl_0,
    g1962_n_spl_
  );


  or

  (
    g1963_n,
    g1940_p_spl_0,
    g1962_p_spl_
  );


  and

  (
    g1964_p,
    g1940_p_spl_,
    g1962_p_spl_
  );


  or

  (
    g1964_n,
    g1940_n_spl_,
    g1962_n_spl_
  );


  and

  (
    g1965_p,
    g1963_n_spl_,
    g1964_n
  );


  or

  (
    g1965_n,
    g1963_p_spl_,
    g1964_p
  );


  and

  (
    g1966_p,
    g1957_n_spl_,
    g1965_p_spl_
  );


  or

  (
    g1966_n,
    g1957_p_spl_,
    g1965_n_spl_
  );


  and

  (
    g1967_p,
    g1957_p_spl_,
    g1965_n_spl_
  );


  or

  (
    g1967_n,
    g1957_n_spl_,
    g1965_p_spl_
  );


  and

  (
    g1968_p,
    g1966_n_spl_,
    g1967_n
  );


  or

  (
    g1968_n,
    g1966_p_spl_,
    g1967_p
  );


  and

  (
    g1969_p,
    g1956_n_spl_,
    g1968_p_spl_
  );


  or

  (
    g1969_n,
    g1956_p_spl_,
    g1968_n_spl_
  );


  and

  (
    g1970_p,
    g1956_p_spl_,
    g1968_n_spl_
  );


  or

  (
    g1970_n,
    g1956_n_spl_,
    g1968_p_spl_
  );


  and

  (
    g1971_p,
    g1969_n_spl_,
    g1970_n
  );


  or

  (
    g1971_n,
    g1969_p_spl_,
    g1970_p
  );


  and

  (
    g1972_p,
    g1955_n_spl_,
    g1971_p_spl_
  );


  or

  (
    g1972_n,
    g1955_p_spl_,
    g1971_n_spl_
  );


  and

  (
    g1973_p,
    g1955_p_spl_,
    g1971_n_spl_
  );


  or

  (
    g1973_n,
    g1955_n_spl_,
    g1971_p_spl_
  );


  and

  (
    g1974_p,
    g1972_n_spl_,
    g1973_n
  );


  or

  (
    g1974_n,
    g1972_p_spl_,
    g1973_p
  );


  or

  (
    g1975_n,
    g1954_p,
    g1974_n
  );


  and

  (
    g1976_p,
    g1969_n_spl_,
    g1972_n_spl_
  );


  or

  (
    g1976_n,
    g1969_p_spl_,
    g1972_p_spl_
  );


  and

  (
    g1977_p,
    G5_p_spl_01,
    G20_p_spl_001
  );


  or

  (
    g1977_n,
    G5_n_spl_1,
    G20_n_spl_001
  );


  and

  (
    g1978_p,
    g1963_n_spl_,
    g1966_n_spl_
  );


  or

  (
    g1978_n,
    g1963_p_spl_,
    g1966_p_spl_
  );


  and

  (
    g1979_p,
    G6_p_spl_01,
    G19_p_spl_010
  );


  or

  (
    g1979_n,
    G6_n_spl_1,
    G19_n_spl_010
  );


  and

  (
    g1980_p,
    G8_p_spl_00,
    G17_p_spl_011
  );


  or

  (
    g1980_n,
    G8_n_spl_0,
    G17_n_spl_011
  );


  and

  (
    g1981_p,
    G7_p_spl_00,
    G18_p_spl_011
  );


  or

  (
    g1981_n,
    G7_n_spl_0,
    G18_n_spl_011
  );


  and

  (
    g1982_p,
    g1980_p_spl_,
    g1981_p_spl_
  );


  or

  (
    g1982_n,
    g1980_n_spl_,
    g1981_n_spl_
  );


  and

  (
    g1983_p,
    g1980_n_spl_,
    g1981_n_spl_
  );


  or

  (
    g1983_n,
    g1980_p_spl_,
    g1981_p_spl_
  );


  and

  (
    g1984_p,
    g1982_n_spl_0,
    g1983_n
  );


  or

  (
    g1984_n,
    g1982_p_spl_0,
    g1983_p
  );


  and

  (
    g1985_p,
    g1960_n_spl_0,
    g1984_n_spl_
  );


  or

  (
    g1985_n,
    g1960_p_spl_0,
    g1984_p_spl_
  );


  and

  (
    g1986_p,
    g1960_p_spl_,
    g1984_p_spl_
  );


  or

  (
    g1986_n,
    g1960_n_spl_,
    g1984_n_spl_
  );


  and

  (
    g1987_p,
    g1985_n_spl_,
    g1986_n
  );


  or

  (
    g1987_n,
    g1985_p_spl_,
    g1986_p
  );


  and

  (
    g1988_p,
    g1979_n_spl_,
    g1987_p_spl_
  );


  or

  (
    g1988_n,
    g1979_p_spl_,
    g1987_n_spl_
  );


  and

  (
    g1989_p,
    g1979_p_spl_,
    g1987_n_spl_
  );


  or

  (
    g1989_n,
    g1979_n_spl_,
    g1987_p_spl_
  );


  and

  (
    g1990_p,
    g1988_n_spl_,
    g1989_n
  );


  or

  (
    g1990_n,
    g1988_p_spl_,
    g1989_p
  );


  and

  (
    g1991_p,
    g1978_n_spl_,
    g1990_p_spl_
  );


  or

  (
    g1991_n,
    g1978_p_spl_,
    g1990_n_spl_
  );


  and

  (
    g1992_p,
    g1978_p_spl_,
    g1990_n_spl_
  );


  or

  (
    g1992_n,
    g1978_n_spl_,
    g1990_p_spl_
  );


  and

  (
    g1993_p,
    g1991_n_spl_,
    g1992_n
  );


  or

  (
    g1993_n,
    g1991_p_spl_,
    g1992_p
  );


  and

  (
    g1994_p,
    g1977_n_spl_,
    g1993_p_spl_
  );


  or

  (
    g1994_n,
    g1977_p_spl_,
    g1993_n_spl_
  );


  and

  (
    g1995_p,
    g1977_p_spl_,
    g1993_n_spl_
  );


  or

  (
    g1995_n,
    g1977_n_spl_,
    g1993_p_spl_
  );


  and

  (
    g1996_p,
    g1994_n_spl_,
    g1995_n
  );


  or

  (
    g1996_n,
    g1994_p_spl_,
    g1995_p
  );


  or

  (
    g1997_n,
    g1976_p,
    g1996_n
  );


  and

  (
    g1998_p,
    g1991_n_spl_,
    g1994_n_spl_
  );


  or

  (
    g1998_n,
    g1991_p_spl_,
    g1994_p_spl_
  );


  and

  (
    g1999_p,
    G6_p_spl_01,
    G20_p_spl_001
  );


  or

  (
    g1999_n,
    G6_n_spl_1,
    G20_n_spl_010
  );


  and

  (
    g2000_p,
    g1985_n_spl_,
    g1988_n_spl_
  );


  or

  (
    g2000_n,
    g1985_p_spl_,
    g1988_p_spl_
  );


  and

  (
    g2001_p,
    G7_p_spl_01,
    G19_p_spl_011
  );


  or

  (
    g2001_n,
    G7_n_spl_1,
    G19_n_spl_011
  );


  and

  (
    g2002_p,
    G9_p_spl_00,
    G17_p_spl_011
  );


  or

  (
    g2002_n,
    G9_n_spl_0,
    G17_n_spl_011
  );


  and

  (
    g2003_p,
    G8_p_spl_00,
    G18_p_spl_011
  );


  or

  (
    g2003_n,
    G8_n_spl_0,
    G18_n_spl_011
  );


  and

  (
    g2004_p,
    g2002_p_spl_,
    g2003_p_spl_
  );


  or

  (
    g2004_n,
    g2002_n_spl_,
    g2003_n_spl_
  );


  and

  (
    g2005_p,
    g2002_n_spl_,
    g2003_n_spl_
  );


  or

  (
    g2005_n,
    g2002_p_spl_,
    g2003_p_spl_
  );


  and

  (
    g2006_p,
    g2004_n_spl_0,
    g2005_n
  );


  or

  (
    g2006_n,
    g2004_p_spl_0,
    g2005_p
  );


  and

  (
    g2007_p,
    g1982_n_spl_0,
    g2006_n_spl_
  );


  or

  (
    g2007_n,
    g1982_p_spl_0,
    g2006_p_spl_
  );


  and

  (
    g2008_p,
    g1982_p_spl_,
    g2006_p_spl_
  );


  or

  (
    g2008_n,
    g1982_n_spl_,
    g2006_n_spl_
  );


  and

  (
    g2009_p,
    g2007_n_spl_,
    g2008_n
  );


  or

  (
    g2009_n,
    g2007_p_spl_,
    g2008_p
  );


  and

  (
    g2010_p,
    g2001_n_spl_,
    g2009_p_spl_
  );


  or

  (
    g2010_n,
    g2001_p_spl_,
    g2009_n_spl_
  );


  and

  (
    g2011_p,
    g2001_p_spl_,
    g2009_n_spl_
  );


  or

  (
    g2011_n,
    g2001_n_spl_,
    g2009_p_spl_
  );


  and

  (
    g2012_p,
    g2010_n_spl_,
    g2011_n
  );


  or

  (
    g2012_n,
    g2010_p_spl_,
    g2011_p
  );


  and

  (
    g2013_p,
    g2000_n_spl_,
    g2012_p_spl_
  );


  or

  (
    g2013_n,
    g2000_p_spl_,
    g2012_n_spl_
  );


  and

  (
    g2014_p,
    g2000_p_spl_,
    g2012_n_spl_
  );


  or

  (
    g2014_n,
    g2000_n_spl_,
    g2012_p_spl_
  );


  and

  (
    g2015_p,
    g2013_n_spl_,
    g2014_n
  );


  or

  (
    g2015_n,
    g2013_p_spl_,
    g2014_p
  );


  and

  (
    g2016_p,
    g1999_n_spl_,
    g2015_p_spl_
  );


  or

  (
    g2016_n,
    g1999_p_spl_,
    g2015_n_spl_
  );


  and

  (
    g2017_p,
    g1999_p_spl_,
    g2015_n_spl_
  );


  or

  (
    g2017_n,
    g1999_n_spl_,
    g2015_p_spl_
  );


  and

  (
    g2018_p,
    g2016_n_spl_,
    g2017_n
  );


  or

  (
    g2018_n,
    g2016_p_spl_,
    g2017_p
  );


  or

  (
    g2019_n,
    g1998_p,
    g2018_n
  );


  and

  (
    g2020_p,
    g2013_n_spl_,
    g2016_n_spl_
  );


  or

  (
    g2020_n,
    g2013_p_spl_,
    g2016_p_spl_
  );


  and

  (
    g2021_p,
    G7_p_spl_01,
    G20_p_spl_010
  );


  or

  (
    g2021_n,
    G7_n_spl_1,
    G20_n_spl_010
  );


  and

  (
    g2022_p,
    g2007_n_spl_,
    g2010_n_spl_
  );


  or

  (
    g2022_n,
    g2007_p_spl_,
    g2010_p_spl_
  );


  and

  (
    g2023_p,
    G8_p_spl_01,
    G19_p_spl_011
  );


  or

  (
    g2023_n,
    G8_n_spl_1,
    G19_n_spl_011
  );


  and

  (
    g2024_p,
    G10_p_spl_00,
    G17_p_spl_100
  );


  or

  (
    g2024_n,
    G10_n_spl_0,
    G17_n_spl_100
  );


  and

  (
    g2025_p,
    G9_p_spl_00,
    G18_p_spl_100
  );


  or

  (
    g2025_n,
    G9_n_spl_0,
    G18_n_spl_100
  );


  and

  (
    g2026_p,
    g2024_p_spl_,
    g2025_p_spl_
  );


  or

  (
    g2026_n,
    g2024_n_spl_,
    g2025_n_spl_
  );


  and

  (
    g2027_p,
    g2024_n_spl_,
    g2025_n_spl_
  );


  or

  (
    g2027_n,
    g2024_p_spl_,
    g2025_p_spl_
  );


  and

  (
    g2028_p,
    g2026_n_spl_0,
    g2027_n
  );


  or

  (
    g2028_n,
    g2026_p_spl_0,
    g2027_p
  );


  and

  (
    g2029_p,
    g2004_n_spl_0,
    g2028_n_spl_
  );


  or

  (
    g2029_n,
    g2004_p_spl_0,
    g2028_p_spl_
  );


  and

  (
    g2030_p,
    g2004_p_spl_,
    g2028_p_spl_
  );


  or

  (
    g2030_n,
    g2004_n_spl_,
    g2028_n_spl_
  );


  and

  (
    g2031_p,
    g2029_n_spl_,
    g2030_n
  );


  or

  (
    g2031_n,
    g2029_p_spl_,
    g2030_p
  );


  and

  (
    g2032_p,
    g2023_n_spl_,
    g2031_p_spl_
  );


  or

  (
    g2032_n,
    g2023_p_spl_,
    g2031_n_spl_
  );


  and

  (
    g2033_p,
    g2023_p_spl_,
    g2031_n_spl_
  );


  or

  (
    g2033_n,
    g2023_n_spl_,
    g2031_p_spl_
  );


  and

  (
    g2034_p,
    g2032_n_spl_,
    g2033_n
  );


  or

  (
    g2034_n,
    g2032_p_spl_,
    g2033_p
  );


  and

  (
    g2035_p,
    g2022_n_spl_,
    g2034_p_spl_
  );


  or

  (
    g2035_n,
    g2022_p_spl_,
    g2034_n_spl_
  );


  and

  (
    g2036_p,
    g2022_p_spl_,
    g2034_n_spl_
  );


  or

  (
    g2036_n,
    g2022_n_spl_,
    g2034_p_spl_
  );


  and

  (
    g2037_p,
    g2035_n_spl_,
    g2036_n
  );


  or

  (
    g2037_n,
    g2035_p_spl_,
    g2036_p
  );


  and

  (
    g2038_p,
    g2021_n_spl_,
    g2037_p_spl_
  );


  or

  (
    g2038_n,
    g2021_p_spl_,
    g2037_n_spl_
  );


  and

  (
    g2039_p,
    g2021_p_spl_,
    g2037_n_spl_
  );


  or

  (
    g2039_n,
    g2021_n_spl_,
    g2037_p_spl_
  );


  and

  (
    g2040_p,
    g2038_n_spl_,
    g2039_n
  );


  or

  (
    g2040_n,
    g2038_p_spl_,
    g2039_p
  );


  or

  (
    g2041_n,
    g2020_p,
    g2040_n
  );


  and

  (
    g2042_p,
    g2035_n_spl_,
    g2038_n_spl_
  );


  or

  (
    g2042_n,
    g2035_p_spl_,
    g2038_p_spl_
  );


  and

  (
    g2043_p,
    G8_p_spl_01,
    G20_p_spl_010
  );


  or

  (
    g2043_n,
    G8_n_spl_1,
    G20_n_spl_011
  );


  and

  (
    g2044_p,
    g2029_n_spl_,
    g2032_n_spl_
  );


  or

  (
    g2044_n,
    g2029_p_spl_,
    g2032_p_spl_
  );


  and

  (
    g2045_p,
    G9_p_spl_01,
    G19_p_spl_100
  );


  or

  (
    g2045_n,
    G9_n_spl_1,
    G19_n_spl_100
  );


  and

  (
    g2046_p,
    G11_p_spl_00,
    G17_p_spl_100
  );


  or

  (
    g2046_n,
    G11_n_spl_0,
    G17_n_spl_100
  );


  and

  (
    g2047_p,
    G10_p_spl_00,
    G18_p_spl_100
  );


  or

  (
    g2047_n,
    G10_n_spl_0,
    G18_n_spl_100
  );


  and

  (
    g2048_p,
    g2046_p_spl_,
    g2047_p_spl_
  );


  or

  (
    g2048_n,
    g2046_n_spl_,
    g2047_n_spl_
  );


  and

  (
    g2049_p,
    g2046_n_spl_,
    g2047_n_spl_
  );


  or

  (
    g2049_n,
    g2046_p_spl_,
    g2047_p_spl_
  );


  and

  (
    g2050_p,
    g2048_n_spl_0,
    g2049_n
  );


  or

  (
    g2050_n,
    g2048_p_spl_0,
    g2049_p
  );


  and

  (
    g2051_p,
    g2026_n_spl_0,
    g2050_n_spl_
  );


  or

  (
    g2051_n,
    g2026_p_spl_0,
    g2050_p_spl_
  );


  and

  (
    g2052_p,
    g2026_p_spl_,
    g2050_p_spl_
  );


  or

  (
    g2052_n,
    g2026_n_spl_,
    g2050_n_spl_
  );


  and

  (
    g2053_p,
    g2051_n_spl_,
    g2052_n
  );


  or

  (
    g2053_n,
    g2051_p_spl_,
    g2052_p
  );


  and

  (
    g2054_p,
    g2045_n_spl_,
    g2053_p_spl_
  );


  or

  (
    g2054_n,
    g2045_p_spl_,
    g2053_n_spl_
  );


  and

  (
    g2055_p,
    g2045_p_spl_,
    g2053_n_spl_
  );


  or

  (
    g2055_n,
    g2045_n_spl_,
    g2053_p_spl_
  );


  and

  (
    g2056_p,
    g2054_n_spl_,
    g2055_n
  );


  or

  (
    g2056_n,
    g2054_p_spl_,
    g2055_p
  );


  and

  (
    g2057_p,
    g2044_n_spl_,
    g2056_p_spl_
  );


  or

  (
    g2057_n,
    g2044_p_spl_,
    g2056_n_spl_
  );


  and

  (
    g2058_p,
    g2044_p_spl_,
    g2056_n_spl_
  );


  or

  (
    g2058_n,
    g2044_n_spl_,
    g2056_p_spl_
  );


  and

  (
    g2059_p,
    g2057_n_spl_,
    g2058_n
  );


  or

  (
    g2059_n,
    g2057_p_spl_,
    g2058_p
  );


  and

  (
    g2060_p,
    g2043_n_spl_,
    g2059_p_spl_
  );


  or

  (
    g2060_n,
    g2043_p_spl_,
    g2059_n_spl_
  );


  and

  (
    g2061_p,
    g2043_p_spl_,
    g2059_n_spl_
  );


  or

  (
    g2061_n,
    g2043_n_spl_,
    g2059_p_spl_
  );


  and

  (
    g2062_p,
    g2060_n_spl_,
    g2061_n
  );


  or

  (
    g2062_n,
    g2060_p_spl_,
    g2061_p
  );


  or

  (
    g2063_n,
    g2042_p,
    g2062_n
  );


  and

  (
    g2064_p,
    g2057_n_spl_,
    g2060_n_spl_
  );


  or

  (
    g2064_n,
    g2057_p_spl_,
    g2060_p_spl_
  );


  and

  (
    g2065_p,
    G9_p_spl_01,
    G20_p_spl_011
  );


  or

  (
    g2065_n,
    G9_n_spl_1,
    G20_n_spl_011
  );


  and

  (
    g2066_p,
    g2051_n_spl_,
    g2054_n_spl_
  );


  or

  (
    g2066_n,
    g2051_p_spl_,
    g2054_p_spl_
  );


  and

  (
    g2067_p,
    G10_p_spl_01,
    G19_p_spl_100
  );


  or

  (
    g2067_n,
    G10_n_spl_1,
    G19_n_spl_100
  );


  and

  (
    g2068_p,
    G12_p_spl_00,
    G17_p_spl_101
  );


  or

  (
    g2068_n,
    G12_n_spl_0,
    G17_n_spl_101
  );


  and

  (
    g2069_p,
    G11_p_spl_00,
    G18_p_spl_101
  );


  or

  (
    g2069_n,
    G11_n_spl_0,
    G18_n_spl_101
  );


  and

  (
    g2070_p,
    g2068_p_spl_,
    g2069_p_spl_
  );


  or

  (
    g2070_n,
    g2068_n_spl_,
    g2069_n_spl_
  );


  and

  (
    g2071_p,
    g2068_n_spl_,
    g2069_n_spl_
  );


  or

  (
    g2071_n,
    g2068_p_spl_,
    g2069_p_spl_
  );


  and

  (
    g2072_p,
    g2070_n_spl_0,
    g2071_n
  );


  or

  (
    g2072_n,
    g2070_p_spl_0,
    g2071_p
  );


  and

  (
    g2073_p,
    g2048_n_spl_0,
    g2072_n_spl_
  );


  or

  (
    g2073_n,
    g2048_p_spl_0,
    g2072_p_spl_
  );


  and

  (
    g2074_p,
    g2048_p_spl_,
    g2072_p_spl_
  );


  or

  (
    g2074_n,
    g2048_n_spl_,
    g2072_n_spl_
  );


  and

  (
    g2075_p,
    g2073_n_spl_,
    g2074_n
  );


  or

  (
    g2075_n,
    g2073_p_spl_,
    g2074_p
  );


  and

  (
    g2076_p,
    g2067_n_spl_,
    g2075_p_spl_
  );


  or

  (
    g2076_n,
    g2067_p_spl_,
    g2075_n_spl_
  );


  and

  (
    g2077_p,
    g2067_p_spl_,
    g2075_n_spl_
  );


  or

  (
    g2077_n,
    g2067_n_spl_,
    g2075_p_spl_
  );


  and

  (
    g2078_p,
    g2076_n_spl_,
    g2077_n
  );


  or

  (
    g2078_n,
    g2076_p_spl_,
    g2077_p
  );


  and

  (
    g2079_p,
    g2066_n_spl_,
    g2078_p_spl_
  );


  or

  (
    g2079_n,
    g2066_p_spl_,
    g2078_n_spl_
  );


  and

  (
    g2080_p,
    g2066_p_spl_,
    g2078_n_spl_
  );


  or

  (
    g2080_n,
    g2066_n_spl_,
    g2078_p_spl_
  );


  and

  (
    g2081_p,
    g2079_n_spl_,
    g2080_n
  );


  or

  (
    g2081_n,
    g2079_p_spl_,
    g2080_p
  );


  and

  (
    g2082_p,
    g2065_n_spl_,
    g2081_p_spl_
  );


  or

  (
    g2082_n,
    g2065_p_spl_,
    g2081_n_spl_
  );


  and

  (
    g2083_p,
    g2065_p_spl_,
    g2081_n_spl_
  );


  or

  (
    g2083_n,
    g2065_n_spl_,
    g2081_p_spl_
  );


  and

  (
    g2084_p,
    g2082_n_spl_,
    g2083_n
  );


  or

  (
    g2084_n,
    g2082_p_spl_,
    g2083_p
  );


  or

  (
    g2085_n,
    g2064_p,
    g2084_n
  );


  and

  (
    g2086_p,
    g2079_n_spl_,
    g2082_n_spl_
  );


  or

  (
    g2086_n,
    g2079_p_spl_,
    g2082_p_spl_
  );


  and

  (
    g2087_p,
    G10_p_spl_01,
    G20_p_spl_011
  );


  or

  (
    g2087_n,
    G10_n_spl_1,
    G20_n_spl_100
  );


  and

  (
    g2088_p,
    g2073_n_spl_,
    g2076_n_spl_
  );


  or

  (
    g2088_n,
    g2073_p_spl_,
    g2076_p_spl_
  );


  and

  (
    g2089_p,
    G11_p_spl_01,
    G19_p_spl_101
  );


  or

  (
    g2089_n,
    G11_n_spl_1,
    G19_n_spl_101
  );


  and

  (
    g2090_p,
    G13_p_spl_00,
    G17_p_spl_101
  );


  or

  (
    g2090_n,
    G13_n_spl_0,
    G17_n_spl_101
  );


  and

  (
    g2091_p,
    G12_p_spl_00,
    G18_p_spl_101
  );


  or

  (
    g2091_n,
    G12_n_spl_0,
    G18_n_spl_101
  );


  and

  (
    g2092_p,
    g2090_p_spl_,
    g2091_p_spl_
  );


  or

  (
    g2092_n,
    g2090_n_spl_,
    g2091_n_spl_
  );


  and

  (
    g2093_p,
    g2090_n_spl_,
    g2091_n_spl_
  );


  or

  (
    g2093_n,
    g2090_p_spl_,
    g2091_p_spl_
  );


  and

  (
    g2094_p,
    g2092_n_spl_0,
    g2093_n
  );


  or

  (
    g2094_n,
    g2092_p_spl_0,
    g2093_p
  );


  and

  (
    g2095_p,
    g2070_n_spl_0,
    g2094_n_spl_
  );


  or

  (
    g2095_n,
    g2070_p_spl_0,
    g2094_p_spl_
  );


  and

  (
    g2096_p,
    g2070_p_spl_,
    g2094_p_spl_
  );


  or

  (
    g2096_n,
    g2070_n_spl_,
    g2094_n_spl_
  );


  and

  (
    g2097_p,
    g2095_n_spl_,
    g2096_n
  );


  or

  (
    g2097_n,
    g2095_p_spl_,
    g2096_p
  );


  and

  (
    g2098_p,
    g2089_n_spl_,
    g2097_p_spl_
  );


  or

  (
    g2098_n,
    g2089_p_spl_,
    g2097_n_spl_
  );


  and

  (
    g2099_p,
    g2089_p_spl_,
    g2097_n_spl_
  );


  or

  (
    g2099_n,
    g2089_n_spl_,
    g2097_p_spl_
  );


  and

  (
    g2100_p,
    g2098_n_spl_,
    g2099_n
  );


  or

  (
    g2100_n,
    g2098_p_spl_,
    g2099_p
  );


  and

  (
    g2101_p,
    g2088_n_spl_,
    g2100_p_spl_
  );


  or

  (
    g2101_n,
    g2088_p_spl_,
    g2100_n_spl_
  );


  and

  (
    g2102_p,
    g2088_p_spl_,
    g2100_n_spl_
  );


  or

  (
    g2102_n,
    g2088_n_spl_,
    g2100_p_spl_
  );


  and

  (
    g2103_p,
    g2101_n_spl_,
    g2102_n
  );


  or

  (
    g2103_n,
    g2101_p_spl_,
    g2102_p
  );


  and

  (
    g2104_p,
    g2087_n_spl_,
    g2103_p_spl_
  );


  or

  (
    g2104_n,
    g2087_p_spl_,
    g2103_n_spl_
  );


  and

  (
    g2105_p,
    g2087_p_spl_,
    g2103_n_spl_
  );


  or

  (
    g2105_n,
    g2087_n_spl_,
    g2103_p_spl_
  );


  and

  (
    g2106_p,
    g2104_n_spl_,
    g2105_n
  );


  or

  (
    g2106_n,
    g2104_p_spl_,
    g2105_p
  );


  or

  (
    g2107_n,
    g2086_p,
    g2106_n
  );


  and

  (
    g2108_p,
    g2101_n_spl_,
    g2104_n_spl_
  );


  or

  (
    g2108_n,
    g2101_p_spl_,
    g2104_p_spl_
  );


  and

  (
    g2109_p,
    G11_p_spl_01,
    G20_p_spl_100
  );


  or

  (
    g2109_n,
    G11_n_spl_1,
    G20_n_spl_100
  );


  and

  (
    g2110_p,
    g2095_n_spl_,
    g2098_n_spl_
  );


  or

  (
    g2110_n,
    g2095_p_spl_,
    g2098_p_spl_
  );


  and

  (
    g2111_p,
    G12_p_spl_01,
    G19_p_spl_101
  );


  or

  (
    g2111_n,
    G12_n_spl_1,
    G19_n_spl_101
  );


  and

  (
    g2112_p,
    G14_p_spl_00,
    G17_p_spl_110
  );


  or

  (
    g2112_n,
    G14_n_spl_0,
    G17_n_spl_110
  );


  and

  (
    g2113_p,
    G13_p_spl_00,
    G18_p_spl_110
  );


  or

  (
    g2113_n,
    G13_n_spl_0,
    G18_n_spl_110
  );


  and

  (
    g2114_p,
    g2112_p_spl_,
    g2113_p_spl_
  );


  or

  (
    g2114_n,
    g2112_n_spl_,
    g2113_n_spl_
  );


  and

  (
    g2115_p,
    g2112_n_spl_,
    g2113_n_spl_
  );


  or

  (
    g2115_n,
    g2112_p_spl_,
    g2113_p_spl_
  );


  and

  (
    g2116_p,
    g2114_n_spl_0,
    g2115_n
  );


  or

  (
    g2116_n,
    g2114_p_spl_0,
    g2115_p
  );


  and

  (
    g2117_p,
    g2092_n_spl_0,
    g2116_n_spl_
  );


  or

  (
    g2117_n,
    g2092_p_spl_0,
    g2116_p_spl_
  );


  and

  (
    g2118_p,
    g2092_p_spl_,
    g2116_p_spl_
  );


  or

  (
    g2118_n,
    g2092_n_spl_,
    g2116_n_spl_
  );


  and

  (
    g2119_p,
    g2117_n_spl_,
    g2118_n
  );


  or

  (
    g2119_n,
    g2117_p_spl_,
    g2118_p
  );


  and

  (
    g2120_p,
    g2111_n_spl_,
    g2119_p_spl_
  );


  or

  (
    g2120_n,
    g2111_p_spl_,
    g2119_n_spl_
  );


  and

  (
    g2121_p,
    g2111_p_spl_,
    g2119_n_spl_
  );


  or

  (
    g2121_n,
    g2111_n_spl_,
    g2119_p_spl_
  );


  and

  (
    g2122_p,
    g2120_n_spl_,
    g2121_n
  );


  or

  (
    g2122_n,
    g2120_p_spl_,
    g2121_p
  );


  and

  (
    g2123_p,
    g2110_n_spl_,
    g2122_p_spl_
  );


  or

  (
    g2123_n,
    g2110_p_spl_,
    g2122_n_spl_
  );


  and

  (
    g2124_p,
    g2110_p_spl_,
    g2122_n_spl_
  );


  or

  (
    g2124_n,
    g2110_n_spl_,
    g2122_p_spl_
  );


  and

  (
    g2125_p,
    g2123_n_spl_,
    g2124_n
  );


  or

  (
    g2125_n,
    g2123_p_spl_,
    g2124_p
  );


  and

  (
    g2126_p,
    g2109_n_spl_,
    g2125_p_spl_
  );


  or

  (
    g2126_n,
    g2109_p_spl_,
    g2125_n_spl_
  );


  and

  (
    g2127_p,
    g2109_p_spl_,
    g2125_n_spl_
  );


  or

  (
    g2127_n,
    g2109_n_spl_,
    g2125_p_spl_
  );


  and

  (
    g2128_p,
    g2126_n_spl_,
    g2127_n
  );


  or

  (
    g2128_n,
    g2126_p_spl_,
    g2127_p
  );


  or

  (
    g2129_n,
    g2108_p,
    g2128_n
  );


  and

  (
    g2130_p,
    g2123_n_spl_,
    g2126_n_spl_
  );


  or

  (
    g2130_n,
    g2123_p_spl_,
    g2126_p_spl_
  );


  and

  (
    g2131_p,
    G12_p_spl_01,
    G20_p_spl_100
  );


  or

  (
    g2131_n,
    G12_n_spl_1,
    G20_n_spl_101
  );


  and

  (
    g2132_p,
    g2117_n_spl_,
    g2120_n_spl_
  );


  or

  (
    g2132_n,
    g2117_p_spl_,
    g2120_p_spl_
  );


  and

  (
    g2133_p,
    G13_p_spl_01,
    G19_p_spl_110
  );


  or

  (
    g2133_n,
    G13_n_spl_1,
    G19_n_spl_110
  );


  and

  (
    g2134_p,
    G15_p_spl_00,
    G17_p_spl_110
  );


  or

  (
    g2134_n,
    G15_n_spl_0,
    G17_n_spl_110
  );


  and

  (
    g2135_p,
    G14_p_spl_00,
    G18_p_spl_110
  );


  or

  (
    g2135_n,
    G14_n_spl_0,
    G18_n_spl_110
  );


  and

  (
    g2136_p,
    g2134_p_spl_,
    g2135_p_spl_
  );


  or

  (
    g2136_n,
    g2134_n_spl_,
    g2135_n_spl_
  );


  and

  (
    g2137_p,
    g2134_n_spl_,
    g2135_n_spl_
  );


  or

  (
    g2137_n,
    g2134_p_spl_,
    g2135_p_spl_
  );


  and

  (
    g2138_p,
    g2136_n_spl_0,
    g2137_n
  );


  or

  (
    g2138_n,
    g2136_p_spl_0,
    g2137_p
  );


  and

  (
    g2139_p,
    g2114_n_spl_0,
    g2138_n_spl_
  );


  or

  (
    g2139_n,
    g2114_p_spl_0,
    g2138_p_spl_
  );


  and

  (
    g2140_p,
    g2114_p_spl_,
    g2138_p_spl_
  );


  or

  (
    g2140_n,
    g2114_n_spl_,
    g2138_n_spl_
  );


  and

  (
    g2141_p,
    g2139_n_spl_,
    g2140_n
  );


  or

  (
    g2141_n,
    g2139_p_spl_,
    g2140_p
  );


  and

  (
    g2142_p,
    g2133_n_spl_,
    g2141_p_spl_
  );


  or

  (
    g2142_n,
    g2133_p_spl_,
    g2141_n_spl_
  );


  and

  (
    g2143_p,
    g2133_p_spl_,
    g2141_n_spl_
  );


  or

  (
    g2143_n,
    g2133_n_spl_,
    g2141_p_spl_
  );


  and

  (
    g2144_p,
    g2142_n_spl_,
    g2143_n
  );


  or

  (
    g2144_n,
    g2142_p_spl_,
    g2143_p
  );


  and

  (
    g2145_p,
    g2132_n_spl_,
    g2144_p_spl_
  );


  or

  (
    g2145_n,
    g2132_p_spl_,
    g2144_n_spl_
  );


  and

  (
    g2146_p,
    g2132_p_spl_,
    g2144_n_spl_
  );


  or

  (
    g2146_n,
    g2132_n_spl_,
    g2144_p_spl_
  );


  and

  (
    g2147_p,
    g2145_n_spl_,
    g2146_n
  );


  or

  (
    g2147_n,
    g2145_p_spl_,
    g2146_p
  );


  and

  (
    g2148_p,
    g2131_n_spl_,
    g2147_p_spl_
  );


  or

  (
    g2148_n,
    g2131_p_spl_,
    g2147_n_spl_
  );


  and

  (
    g2149_p,
    g2131_p_spl_,
    g2147_n_spl_
  );


  or

  (
    g2149_n,
    g2131_n_spl_,
    g2147_p_spl_
  );


  and

  (
    g2150_p,
    g2148_n_spl_,
    g2149_n
  );


  or

  (
    g2150_n,
    g2148_p_spl_,
    g2149_p
  );


  or

  (
    g2151_n,
    g2130_p,
    g2150_n
  );


  and

  (
    g2152_p,
    g2145_n_spl_,
    g2148_n_spl_
  );


  or

  (
    g2152_n,
    g2145_p_spl_,
    g2148_p_spl_
  );


  and

  (
    g2153_p,
    G13_p_spl_01,
    G20_p_spl_101
  );


  or

  (
    g2153_n,
    G13_n_spl_1,
    G20_n_spl_101
  );


  and

  (
    g2154_p,
    g2139_n_spl_,
    g2142_n_spl_
  );


  or

  (
    g2154_n,
    g2139_p_spl_,
    g2142_p_spl_
  );


  and

  (
    g2155_p,
    G14_p_spl_01,
    G19_p_spl_110
  );


  or

  (
    g2155_n,
    G14_n_spl_1,
    G19_n_spl_110
  );


  and

  (
    g2156_p,
    G16_p_spl_00,
    G17_p_spl_111
  );


  or

  (
    g2156_n,
    G16_n_spl_0,
    G17_n_spl_11
  );


  and

  (
    g2157_p,
    G15_p_spl_00,
    G18_p_spl_111
  );


  or

  (
    g2157_n,
    G15_n_spl_0,
    G18_n_spl_111
  );


  and

  (
    g2158_p,
    g2156_p_spl_,
    g2157_p_spl_
  );


  or

  (
    g2158_n,
    g2156_n_spl_,
    g2157_n_spl_
  );


  and

  (
    g2159_p,
    g2156_n_spl_,
    g2157_n_spl_
  );


  or

  (
    g2159_n,
    g2156_p_spl_,
    g2157_p_spl_
  );


  and

  (
    g2160_p,
    g2158_n_spl_,
    g2159_n
  );


  or

  (
    g2160_n,
    g2158_p_spl_,
    g2159_p
  );


  and

  (
    g2161_p,
    g2136_n_spl_0,
    g2160_n_spl_
  );


  or

  (
    g2161_n,
    g2136_p_spl_0,
    g2160_p_spl_
  );


  and

  (
    g2162_p,
    g2136_p_spl_,
    g2160_p_spl_
  );


  or

  (
    g2162_n,
    g2136_n_spl_,
    g2160_n_spl_
  );


  and

  (
    g2163_p,
    g2161_n_spl_,
    g2162_n
  );


  or

  (
    g2163_n,
    g2161_p_spl_,
    g2162_p
  );


  and

  (
    g2164_p,
    g2155_n_spl_,
    g2163_p_spl_
  );


  or

  (
    g2164_n,
    g2155_p_spl_,
    g2163_n_spl_
  );


  and

  (
    g2165_p,
    g2155_p_spl_,
    g2163_n_spl_
  );


  or

  (
    g2165_n,
    g2155_n_spl_,
    g2163_p_spl_
  );


  and

  (
    g2166_p,
    g2164_n_spl_,
    g2165_n
  );


  or

  (
    g2166_n,
    g2164_p_spl_,
    g2165_p
  );


  and

  (
    g2167_p,
    g2154_n_spl_,
    g2166_p_spl_
  );


  or

  (
    g2167_n,
    g2154_p_spl_,
    g2166_n_spl_
  );


  and

  (
    g2168_p,
    g2154_p_spl_,
    g2166_n_spl_
  );


  or

  (
    g2168_n,
    g2154_n_spl_,
    g2166_p_spl_
  );


  and

  (
    g2169_p,
    g2167_n_spl_,
    g2168_n
  );


  or

  (
    g2169_n,
    g2167_p_spl_,
    g2168_p
  );


  and

  (
    g2170_p,
    g2153_n_spl_,
    g2169_p_spl_
  );


  or

  (
    g2170_n,
    g2153_p_spl_,
    g2169_n_spl_
  );


  and

  (
    g2171_p,
    g2153_p_spl_,
    g2169_n_spl_
  );


  or

  (
    g2171_n,
    g2153_n_spl_,
    g2169_p_spl_
  );


  and

  (
    g2172_p,
    g2170_n_spl_,
    g2171_n
  );


  or

  (
    g2172_n,
    g2170_p_spl_,
    g2171_p
  );


  or

  (
    g2173_n,
    g2152_p,
    g2172_n
  );


  and

  (
    g2174_p,
    g2167_n_spl_,
    g2170_n_spl_
  );


  or

  (
    g2174_n,
    g2167_p_spl_,
    g2170_p_spl_
  );


  and

  (
    g2175_p,
    G14_p_spl_01,
    G20_p_spl_101
  );


  or

  (
    g2175_n,
    G14_n_spl_1,
    G20_n_spl_110
  );


  and

  (
    g2176_p,
    g2161_n_spl_,
    g2164_n_spl_
  );


  or

  (
    g2176_n,
    g2161_p_spl_,
    g2164_p_spl_
  );


  and

  (
    g2177_p,
    G16_p_spl_00,
    G18_p_spl_111
  );


  or

  (
    g2177_n,
    G16_n_spl_0,
    G18_n_spl_111
  );


  and

  (
    g2178_p,
    g2158_n_spl_,
    g2177_p_spl_
  );


  or

  (
    g2178_n,
    g2158_p_spl_,
    g2177_n_spl_
  );


  and

  (
    g2179_p,
    G15_p_spl_0,
    G19_p_spl_111
  );


  or

  (
    g2179_n,
    G15_n_spl_1,
    G19_n_spl_111
  );


  and

  (
    g2180_p,
    g2178_p_spl_,
    g2179_n_spl_
  );


  or

  (
    g2180_n,
    g2178_n_spl_,
    g2179_p_spl_
  );


  and

  (
    g2181_p,
    g2178_n_spl_,
    g2179_p_spl_
  );


  or

  (
    g2181_n,
    g2178_p_spl_,
    g2179_n_spl_
  );


  and

  (
    g2182_p,
    g2180_n_spl_,
    g2181_n
  );


  or

  (
    g2182_n,
    g2180_p_spl_,
    g2181_p
  );


  and

  (
    g2183_p,
    g2176_n_spl_,
    g2182_p_spl_
  );


  or

  (
    g2183_n,
    g2176_p_spl_,
    g2182_n_spl_
  );


  and

  (
    g2184_p,
    g2176_p_spl_,
    g2182_n_spl_
  );


  or

  (
    g2184_n,
    g2176_n_spl_,
    g2182_p_spl_
  );


  and

  (
    g2185_p,
    g2183_n_spl_,
    g2184_n
  );


  or

  (
    g2185_n,
    g2183_p_spl_,
    g2184_p
  );


  and

  (
    g2186_p,
    g2175_n_spl_,
    g2185_p_spl_
  );


  or

  (
    g2186_n,
    g2175_p_spl_,
    g2185_n_spl_
  );


  and

  (
    g2187_p,
    g2175_p_spl_,
    g2185_n_spl_
  );


  or

  (
    g2187_n,
    g2175_n_spl_,
    g2185_p_spl_
  );


  and

  (
    g2188_p,
    g2186_n_spl_,
    g2187_n
  );


  or

  (
    g2188_n,
    g2186_p_spl_,
    g2187_p
  );


  or

  (
    g2189_n,
    g2174_p,
    g2188_n
  );


  and

  (
    g2190_p,
    g2183_n_spl_,
    g2186_n_spl_
  );


  or

  (
    g2190_n,
    g2183_p_spl_,
    g2186_p_spl_
  );


  and

  (
    g2191_p,
    G15_p_spl_1,
    G20_p_spl_110
  );


  or

  (
    g2191_n,
    G15_n_spl_1,
    G20_n_spl_110
  );


  and

  (
    g2192_p,
    G16_p_spl_0,
    G19_p_spl_111
  );


  or

  (
    g2192_n,
    G16_n_spl_,
    G19_n_spl_111
  );


  and

  (
    g2193_p,
    g2177_p_spl_,
    g2180_n_spl_
  );


  or

  (
    g2193_n,
    g2177_n_spl_,
    g2180_p_spl_
  );


  and

  (
    g2194_p,
    g2192_n_spl_,
    g2193_n_spl_
  );


  or

  (
    g2194_n,
    g2192_p_spl_,
    g2193_p_spl_
  );


  and

  (
    g2195_p,
    g2192_p_spl_,
    g2193_p_spl_
  );


  or

  (
    g2195_n,
    g2192_n_spl_,
    g2193_n_spl_
  );


  and

  (
    g2196_p,
    g2194_n_spl_,
    g2195_n
  );


  or

  (
    g2196_n,
    g2194_p,
    g2195_p
  );


  and

  (
    g2197_p,
    g2191_n_spl_,
    g2196_p_spl_
  );


  or

  (
    g2197_n,
    g2191_p_spl_,
    g2196_n_spl_
  );


  and

  (
    g2198_p,
    g2191_p_spl_,
    g2196_n_spl_
  );


  or

  (
    g2198_n,
    g2191_n_spl_,
    g2196_p_spl_
  );


  and

  (
    g2199_p,
    g2197_n_spl_,
    g2198_n
  );


  or

  (
    g2199_n,
    g2197_p,
    g2198_p
  );


  or

  (
    g2200_n,
    g2190_p,
    g2199_n
  );


  and

  (
    g2201_p,
    g1585_n_spl_,
    g1588_n_spl_
  );


  or

  (
    g2201_n,
    g1585_p_spl_,
    g1588_p_spl_
  );


  and

  (
    g2202_p,
    g1932_p_spl_,
    g1934_n_spl_
  );


  or

  (
    g2202_n,
    g1932_n_spl_,
    g1934_p_spl_
  );


  and

  (
    g2203_p,
    g1935_n_spl_,
    g2202_n
  );


  or

  (
    g2203_n,
    g1935_p_spl_,
    g2202_p
  );


  and

  (
    g2204_p,
    g2201_n_spl_,
    g2203_p_spl_
  );


  or

  (
    g2204_n,
    g2201_p_spl_,
    g2203_n_spl_
  );


  and

  (
    g2205_p,
    G2_p_spl_01,
    G20_p_spl_110
  );


  or

  (
    g2205_n,
    G2_n_spl_1,
    G20_n_spl_11
  );


  and

  (
    g2206_p,
    g2201_p_spl_,
    g2203_n_spl_
  );


  or

  (
    g2206_n,
    g2201_n_spl_,
    g2203_p_spl_
  );


  and

  (
    g2207_p,
    g2204_n_spl_,
    g2206_n
  );


  or

  (
    g2207_n,
    g2204_p_spl_,
    g2206_p
  );


  and

  (
    g2208_p,
    g2205_n_spl_,
    g2207_p_spl_
  );


  or

  (
    g2208_n,
    g2205_p,
    g2207_n
  );


  and

  (
    g2209_p,
    g2204_n_spl_,
    g2208_n_spl_
  );


  or

  (
    g2209_n,
    g2204_p_spl_,
    g2208_p
  );


  and

  (
    g2210_p,
    g1950_p_spl_,
    g1952_n_spl_
  );


  or

  (
    g2210_n,
    g1950_n_spl_,
    g1952_p_spl_
  );


  and

  (
    g2211_p,
    g1953_n_spl_,
    g2210_n
  );


  or

  (
    g2211_n,
    g1953_p_spl_,
    g2210_p
  );


  or

  (
    g2212_n,
    g2209_p,
    g2211_n
  );


  and

  (
    g2213_p,
    G3_p_spl_1,
    G21_p_spl_000
  );


  and

  (
    g2214_p,
    G4_p_spl_1,
    G21_p_spl_000
  );


  and

  (
    g2215_p,
    G5_p_spl_1,
    G21_p_spl_001
  );


  and

  (
    g2216_p,
    G6_p_spl_1,
    G21_p_spl_001
  );


  and

  (
    g2217_p,
    G7_p_spl_1,
    G21_p_spl_010
  );


  and

  (
    g2218_p,
    G8_p_spl_1,
    G21_p_spl_010
  );


  and

  (
    g2219_p,
    G9_p_spl_1,
    G21_p_spl_011
  );


  and

  (
    g2220_p,
    G10_p_spl_1,
    G21_p_spl_011
  );


  and

  (
    g2221_p,
    G11_p_spl_1,
    G21_p_spl_100
  );


  and

  (
    g2222_p,
    G12_p_spl_1,
    G21_p_spl_100
  );


  and

  (
    g2223_p,
    G13_p_spl_1,
    G21_p_spl_101
  );


  and

  (
    g2224_p,
    G14_p_spl_1,
    G21_p_spl_101
  );


  and

  (
    g2225_p,
    G16_p_spl_1,
    G20_p_spl_11
  );


  and

  (
    g2226_p,
    G2_p_spl_1,
    G21_p_spl_11
  );


  and

  (
    g2227_p,
    g2194_n_spl_,
    g2197_n_spl_
  );


  or

  (
    g2228_n,
    g1591_p,
    g1631_p_spl_
  );


  or

  (
    g2229_n,
    g2205_n_spl_,
    g2207_p_spl_
  );


  and

  (
    g2230_p,
    g2208_n_spl_,
    g2229_n
  );


  and

  (
    g2231_p,
    g2228_n_spl_,
    g2230_p_spl_
  );


  or

  (
    g2232_n,
    g2228_n_spl_,
    g2230_p_spl_
  );


  or

  (
    g2233_n,
    g1954_n,
    g1974_p
  );


  and

  (
    g2234_p,
    g1975_n_spl_,
    g2233_n
  );


  or

  (
    g2235_n,
    g1976_n,
    g1996_p
  );


  and

  (
    g2236_p,
    g1997_n_spl_,
    g2235_n
  );


  or

  (
    g2237_n,
    g1998_n,
    g2018_p
  );


  and

  (
    g2238_p,
    g2019_n_spl_,
    g2237_n
  );


  or

  (
    g2239_n,
    g2020_n,
    g2040_p
  );


  and

  (
    g2240_p,
    g2041_n_spl_,
    g2239_n
  );


  or

  (
    g2241_n,
    g2042_n,
    g2062_p
  );


  and

  (
    g2242_p,
    g2063_n_spl_,
    g2241_n
  );


  or

  (
    g2243_n,
    g2064_n,
    g2084_p
  );


  and

  (
    g2244_p,
    g2085_n_spl_,
    g2243_n
  );


  or

  (
    g2245_n,
    g2086_n,
    g2106_p
  );


  and

  (
    g2246_p,
    g2107_n_spl_,
    g2245_n
  );


  or

  (
    g2247_n,
    g2108_n,
    g2128_p
  );


  and

  (
    g2248_p,
    g2129_n_spl_,
    g2247_n
  );


  or

  (
    g2249_n,
    g2130_n,
    g2150_p
  );


  and

  (
    g2250_p,
    g2151_n_spl_,
    g2249_n
  );


  or

  (
    g2251_n,
    g2152_n,
    g2172_p
  );


  and

  (
    g2252_p,
    g2173_n_spl_,
    g2251_n
  );


  or

  (
    g2253_n,
    g2174_n,
    g2188_p
  );


  and

  (
    g2254_p,
    g2189_n_spl_,
    g2253_n
  );


  or

  (
    g2255_n,
    g2190_n,
    g2199_p
  );


  and

  (
    g2256_p,
    g2200_n_spl_,
    g2255_n
  );


  or

  (
    g2257_n,
    g2209_n,
    g2211_p
  );


  and

  (
    g2258_p,
    g2212_n_spl_,
    g2257_n
  );


  buf

  (
    G6257,
    g389_p
  );


  buf

  (
    G6258,
    g391_p
  );


  buf

  (
    G6259,
    g393_n
  );


  buf

  (
    G6260,
    g395_n
  );


  buf

  (
    G6261,
    g397_n
  );


  buf

  (
    G6262,
    g399_n
  );


  buf

  (
    G6263,
    g401_n
  );


  buf

  (
    G6264,
    g403_n
  );


  buf

  (
    G6265,
    g405_n
  );


  buf

  (
    G6266,
    g407_n
  );


  buf

  (
    G6267,
    g409_n
  );


  buf

  (
    G6268,
    g411_n
  );


  buf

  (
    G6269,
    g413_n
  );


  buf

  (
    G6270,
    g415_n
  );


  buf

  (
    G6271,
    g417_n
  );


  buf

  (
    G6272,
    g419_n
  );


  buf

  (
    G6273,
    g421_p
  );


  buf

  (
    G6274,
    g423_n
  );


  buf

  (
    G6275,
    g425_n
  );


  buf

  (
    G6276,
    g427_n
  );


  buf

  (
    G6277,
    g429_n
  );


  buf

  (
    G6278,
    g431_n
  );


  buf

  (
    G6279,
    g436_n
  );


  buf

  (
    G6280,
    g445_n
  );


  buf

  (
    G6281,
    g458_n
  );


  buf

  (
    G6282,
    g475_n
  );


  buf

  (
    G6283,
    g496_n
  );


  buf

  (
    G6284,
    g521_n
  );


  buf

  (
    G6285,
    g546_n
  );


  buf

  (
    G6286,
    g563_n
  );


  buf

  (
    G6287,
    g571_p
  );


  not

  (
    G6288,
    g573_p
  );


  buf

  (
    n5322_li003_li003,
    n4908_o2_p_spl_
  );


  buf

  (
    n5430_li039_li039,
    n4843_o2_p_spl_1
  );


  buf

  (
    n5442_li043_li043,
    n4844_o2_p_spl_1
  );


  buf

  (
    n5454_li047_li047,
    n4845_o2_p_spl_
  );


  buf

  (
    n5466_li051_li051,
    n4846_o2_p_spl_1
  );


  buf

  (
    n5478_li055_li055,
    n4847_o2_p_spl_1
  );


  buf

  (
    n5490_li059_li059,
    n4848_o2_p_spl_
  );


  buf

  (
    n5502_li063_li063,
    n4849_o2_p_spl_1
  );


  buf

  (
    n5514_li067_li067,
    n4850_o2_p
  );


  buf

  (
    n5565_li084_li084,
    G22_p
  );


  buf

  (
    n5577_li088_li088,
    G23_p
  );


  buf

  (
    n5589_li092_li092,
    G24_p
  );


  buf

  (
    n5601_li096_li096,
    G25_p
  );


  buf

  (
    n5613_li100_li100,
    G26_p
  );


  buf

  (
    n5625_li104_li104,
    G27_p
  );


  buf

  (
    n5628_li105_li105,
    n2794_lo_p
  );


  buf

  (
    n5637_li108_li108,
    G28_p
  );


  buf

  (
    n5640_li109_li109,
    n2806_lo_p
  );


  buf

  (
    n5649_li112_li112,
    G29_p
  );


  buf

  (
    n5652_li113_li113,
    n2818_lo_p
  );


  buf

  (
    n5661_li116_li116,
    G30_p
  );


  buf

  (
    n5664_li117_li117,
    n2830_lo_p
  );


  buf

  (
    n5670_li119_li119,
    lo118_buf_o2_p_spl_11
  );


  buf

  (
    n5673_li120_li120,
    G31_p
  );


  buf

  (
    n5676_li121_li121,
    n2842_lo_p
  );


  buf

  (
    n5679_li122_li122,
    n2845_lo_p
  );


  buf

  (
    n5682_li123_li123,
    n2848_lo_p_spl_11
  );


  buf

  (
    n5685_li124_li124,
    G32_p
  );


  buf

  (
    n5688_li125_li125,
    n2854_lo_p
  );


  buf

  (
    n5691_li126_li126,
    n2857_lo_p
  );


  buf

  (
    n5694_li127_li127,
    n2860_lo_p_spl_11
  );


  buf

  (
    n3737_i2,
    n4960_o2_p
  );


  buf

  (
    n3736_i2,
    n316_inv_p
  );


  buf

  (
    n3801_i2,
    n325_inv_p
  );


  buf

  (
    n3836_i2,
    n328_inv_p
  );


  buf

  (
    n3885_i2,
    n331_inv_p
  );


  buf

  (
    n3902_i2,
    n5189_o2_p
  );


  buf

  (
    n4002_i2,
    n340_inv_p
  );


  buf

  (
    n4052_i2,
    n346_inv_p
  );


  buf

  (
    n4067_i2,
    n5388_o2_p
  );


  buf

  (
    n4162_i2,
    n355_inv_p
  );


  buf

  (
    n4212_i2,
    n358_inv_p
  );


  buf

  (
    n4227_i2,
    n5612_o2_p
  );


  buf

  (
    n4321_i2,
    n367_inv_p
  );


  buf

  (
    n4367_i2,
    n373_inv_p
  );


  buf

  (
    n4383_i2,
    n5802_o2_p
  );


  buf

  (
    n4475_i2,
    n382_inv_p
  );


  buf

  (
    n4523_i2,
    n385_inv_p
  );


  buf

  (
    n4537_i2,
    n6023_o2_p
  );


  buf

  (
    n4628_i2,
    n394_inv_p
  );


  buf

  (
    n4674_i2,
    n400_inv_p
  );


  buf

  (
    n4688_i2,
    n6383_o2_p
  );


  buf

  (
    n4791_i2,
    n409_inv_p
  );


  buf

  (
    n4835_i2,
    n418_inv_p
  );


  buf

  (
    n4868_i2,
    n6726_o2_p
  );


  buf

  (
    n5086_i2,
    n490_inv_p
  );


  buf

  (
    n5130_i2,
    n499_inv_p
  );


  buf

  (
    n5188_i2,
    n772_o2_p
  );


  buf

  (
    n5402_i2,
    n529_inv_p
  );


  buf

  (
    n5445_i2,
    n535_inv_p
  );


  buf

  (
    n5500_i2,
    n848_o2_p
  );


  buf

  (
    n5707_i2,
    n559_inv_p
  );


  buf

  (
    n5745_i2,
    n577_inv_p
  );


  buf

  (
    n5801_i2,
    n932_o2_p
  );


  buf

  (
    n4836_i2,
    n6024_o2_p_spl_1
  );


  buf

  (
    n4837_i2,
    n6025_o2_p_spl_1
  );


  buf

  (
    n4838_i2,
    n6026_o2_p_spl_1
  );


  buf

  (
    n4839_i2,
    n6027_o2_p_spl_1
  );


  buf

  (
    n4840_i2,
    n6028_o2_p_spl_1
  );


  buf

  (
    n4841_i2,
    n6029_o2_p_spl_1
  );


  buf

  (
    n4842_i2,
    n6030_o2_p_spl_1
  );


  buf

  (
    n4843_i2,
    n6031_o2_p_spl_1
  );


  buf

  (
    n4844_i2,
    n6032_o2_p_spl_1
  );


  buf

  (
    n4845_i2,
    n6033_o2_p_spl_1
  );


  buf

  (
    n4846_i2,
    n6034_o2_p_spl_1
  );


  buf

  (
    n4847_i2,
    n6035_o2_p_spl_1
  );


  buf

  (
    n4848_i2,
    n6036_o2_p_spl_1
  );


  buf

  (
    n4849_i2,
    n6037_o2_p_spl_1
  );


  buf

  (
    n4850_i2,
    n6038_o2_p
  );


  buf

  (
    n4867_i2,
    n6053_o2_p_spl_1
  );


  buf

  (
    n4908_i2,
    n6148_o2_p_spl_1
  );


  buf

  (
    n6081_i2,
    n655_inv_p
  );


  buf

  (
    n6120_i2,
    n682_inv_p
  );


  buf

  (
    n4959_i2,
    n481_inv_p
  );


  buf

  (
    n4960_i2,
    n6201_o2_p
  );


  buf

  (
    n6203_i2,
    n1024_o2_p
  );


  buf

  (
    n5040_i2,
    n487_inv_p
  );


  buf

  (
    n5087_i2,
    n493_inv_p
  );


  buf

  (
    n5158_i2,
    n502_inv_p
  );


  buf

  (
    n5189_i2,
    n6482_o2_p
  );


  buf

  (
    n6594_i2,
    n754_inv_p
  );


  buf

  (
    n5328_i2,
    n520_inv_p
  );


  buf

  (
    n6631_i2,
    n829_inv_p
  );


  buf

  (
    n5372_i2,
    n523_inv_p
  );


  buf

  (
    n5388_i2,
    n6727_o2_p
  );


  buf

  (
    n6725_i2,
    n1124_o2_p_spl_
  );


  buf

  (
    n5527_i2,
    n541_inv_p
  );


  buf

  (
    n5555_i2,
    n544_inv_p
  );


  buf

  (
    n5612_i2,
    n512_o2_p
  );


  buf

  (
    n1127_i2,
    g574_p_spl_
  );


  buf

  (
    n5708_i2,
    n562_inv_p
  );


  buf

  (
    n1231_i2,
    g579_p_spl_
  );


  buf

  (
    n5771_i2,
    n580_inv_p
  );


  buf

  (
    n5802_i2,
    n548_o2_p
  );


  buf

  (
    n1232_i2,
    g580_p_spl_
  );


  buf

  (
    n5948_i2,
    n598_inv_p
  );


  buf

  (
    n6006_i2,
    n601_inv_p
  );


  buf

  (
    n6023_i2,
    n592_o2_p
  );


  not

  (
    n1235_i2,
    g581_n_spl_
  );


  buf

  (
    n6243_i2,
    n700_inv_p
  );


  buf

  (
    n1347_i2,
    g592_p_spl_
  );


  buf

  (
    n6296_i2,
    n706_inv_p
  );


  buf

  (
    n6383_i2,
    n644_o2_p
  );


  buf

  (
    n1348_i2,
    g593_p_spl_
  );


  buf

  (
    n6595_i2,
    n757_inv_p
  );


  not

  (
    n1351_i2,
    g594_n_spl_
  );


  not

  (
    n1461_i2,
    g609_p_spl_
  );


  buf

  (
    n6655_i2,
    n844_inv_p
  );


  buf

  (
    n6024_i2,
    lo010_buf_o2_p_spl_1
  );


  buf

  (
    n6025_i2,
    lo014_buf_o2_p_spl_1
  );


  buf

  (
    n6026_i2,
    lo018_buf_o2_p_spl_1
  );


  buf

  (
    n6027_i2,
    lo022_buf_o2_p_spl_1
  );


  buf

  (
    n6028_i2,
    lo026_buf_o2_p_spl_1
  );


  buf

  (
    n6029_i2,
    lo030_buf_o2_p_spl_1
  );


  buf

  (
    n6030_i2,
    lo034_buf_o2_p_spl_1
  );


  buf

  (
    n6031_i2,
    lo038_buf_o2_p_spl_1
  );


  buf

  (
    n6032_i2,
    lo042_buf_o2_p_spl_1
  );


  buf

  (
    n6033_i2,
    lo046_buf_o2_p_spl_1
  );


  buf

  (
    n6034_i2,
    lo050_buf_o2_p_spl_1
  );


  buf

  (
    n6035_i2,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    n6036_i2,
    lo058_buf_o2_p_spl_1
  );


  buf

  (
    n6037_i2,
    lo062_buf_o2_p_spl_
  );


  buf

  (
    n6038_i2,
    lo066_buf_o2_p
  );


  buf

  (
    n6053_i2,
    lo006_buf_o2_p_spl_1
  );


  buf

  (
    n6726_i2,
    n704_o2_p
  );


  buf

  (
    n6148_i2,
    lo002_buf_o2_p_spl_1
  );


  not

  (
    n1463_i2,
    g610_n_spl_
  );


  buf

  (
    n1573_i2,
    g629_p_spl_
  );


  buf

  (
    n6200_i2,
    n691_inv_p
  );


  buf

  (
    n6201_i2,
    n451_o2_p
  );


  buf

  (
    n6294_i2,
    n703_inv_p
  );


  buf

  (
    n707_i2,
    g630_p_spl_
  );


  buf

  (
    n6361_i2,
    n718_inv_p
  );


  buf

  (
    n1574_i2,
    g631_p_spl_
  );


  buf

  (
    n771_i2,
    g634_p_spl_
  );


  buf

  (
    n6423_i2,
    n736_inv_p
  );


  buf

  (
    n772_i2,
    g635_p_spl_
  );


  buf

  (
    n6482_i2,
    n464_o2_p
  );


  buf

  (
    lo106_buf_i2,
    n2797_lo_p_spl_111
  );


  not

  (
    n1577_i2,
    g636_n_spl_
  );


  buf

  (
    n1678_i2,
    g659_p_spl_
  );


  buf

  (
    n6596_i2,
    n760_inv_p
  );


  buf

  (
    n6683_i2,
    n847_inv_p
  );


  buf

  (
    n6727_i2,
    n484_o2_p
  );


  buf

  (
    n775_i2,
    g660_p_spl_
  );


  buf

  (
    n1679_i2,
    g661_p_spl_
  );


  buf

  (
    n847_i2,
    g670_p_spl_
  );


  buf

  (
    n848_i2,
    g671_p_spl_
  );


  buf

  (
    n487_i2,
    g672_p_spl_
  );


  buf

  (
    n511_i2,
    g673_p_spl_
  );


  buf

  (
    lo110_buf_i2,
    n2809_lo_p_spl_11
  );


  not

  (
    n1682_i2,
    g674_n_spl_
  );


  buf

  (
    n1775_i2,
    g701_p_spl_
  );


  buf

  (
    n512_i2,
    g702_p_spl_
  );


  buf

  (
    n851_i2,
    g703_p_spl_
  );


  buf

  (
    n515_i2,
    g704_p_spl_
  );


  buf

  (
    n2210_i2,
    g739_n_spl_
  );


  buf

  (
    n2126_i2,
    g789_n_spl_
  );


  buf

  (
    n2010_i2,
    g839_n_spl_
  );


  buf

  (
    n1776_i2,
    g840_p_spl_
  );


  buf

  (
    n931_i2,
    g857_p_spl_
  );


  buf

  (
    n547_i2,
    g864_p_spl_
  );


  buf

  (
    n932_i2,
    g865_p_spl_
  );


  buf

  (
    n548_i2,
    g866_p_spl_
  );


  buf

  (
    lo114_buf_i2,
    n2821_lo_p_spl_11
  );


  not

  (
    n1779_i2,
    g867_n_spl_
  );


  buf

  (
    n1864_i2,
    g889_p_spl_
  );


  buf

  (
    n551_i2,
    g890_p_spl_
  );


  buf

  (
    n591_i2,
    g905_p_spl_
  );


  buf

  (
    n592_i2,
    g906_p_spl_
  );


  buf

  (
    lo010_buf_i2,
    G3_p_spl_1
  );


  buf

  (
    lo014_buf_i2,
    G4_p_spl_1
  );


  buf

  (
    lo018_buf_i2,
    G5_p_spl_1
  );


  buf

  (
    lo022_buf_i2,
    G6_p_spl_1
  );


  buf

  (
    lo026_buf_i2,
    G7_p_spl_1
  );


  buf

  (
    lo030_buf_i2,
    G8_p_spl_1
  );


  buf

  (
    lo034_buf_i2,
    G9_p_spl_1
  );


  buf

  (
    lo038_buf_i2,
    G10_p_spl_1
  );


  buf

  (
    lo042_buf_i2,
    G11_p_spl_1
  );


  buf

  (
    lo046_buf_i2,
    G12_p_spl_1
  );


  buf

  (
    lo050_buf_i2,
    G13_p_spl_1
  );


  buf

  (
    lo054_buf_i2,
    G14_p_spl_1
  );


  buf

  (
    lo058_buf_i2,
    G15_p_spl_1
  );


  buf

  (
    lo062_buf_i2,
    G16_p_spl_1
  );


  buf

  (
    lo066_buf_i2,
    G17_p_spl_111
  );


  buf

  (
    lo006_buf_i2,
    G2_p_spl_1
  );


  buf

  (
    n935_i2,
    g907_p_spl_
  );


  not

  (
    n2013_i2,
    g911_n_spl_
  );


  not

  (
    n2129_i2,
    g915_n_spl_
  );


  not

  (
    n2213_i2,
    g919_n_spl_
  );


  buf

  (
    n2243_i2,
    g922_n_spl_
  );


  buf

  (
    n2175_i2,
    g934_n_spl_
  );


  buf

  (
    n2075_i2,
    g946_n_spl_
  );


  buf

  (
    n1943_i2,
    g958_n_spl_
  );


  buf

  (
    n1865_i2,
    g959_p_spl_
  );


  buf

  (
    n1023_i2,
    g984_p_spl_
  );


  buf

  (
    lo094_buf_i2,
    n2758_lo_p_spl_11
  );


  buf

  (
    lo002_buf_i2,
    G1_p_spl_
  );


  buf

  (
    n450_i2,
    g985_p_spl_
  );


  buf

  (
    n451_i2,
    g986_p_spl_
  );


  buf

  (
    n1024_i2,
    g987_p_spl_
  );


  buf

  (
    n595_i2,
    g988_p_spl_
  );


  buf

  (
    n452_i2,
    g989_p_spl_
  );


  buf

  (
    n643_i2,
    g1012_p_spl_
  );


  buf

  (
    lo118_buf_i2,
    n2833_lo_p_spl_1
  );


  not

  (
    n1868_i2,
    g1013_n_spl_
  );


  buf

  (
    n1945_i2,
    g1015_p_spl_
  );


  buf

  (
    n455_i2,
    g1016_p_spl_
  );


  buf

  (
    n2045_i2,
    g1053_n_spl_
  );


  buf

  (
    n1913_i2,
    g1107_n_spl_
  );


  buf

  (
    n1749_i2,
    g1164_n_spl_
  );


  buf

  (
    n1553_i2,
    g1241_n_spl_
  );


  buf

  (
    n644_i2,
    g1242_p_spl_
  );


  buf

  (
    n463_i2,
    g1250_p_spl_
  );


  buf

  (
    lo098_buf_i2,
    n2770_lo_p_spl_11
  );


  buf

  (
    n1121_i2,
    g1278_n_spl_
  );


  buf

  (
    n1719_i2,
    g1328_n_spl_
  );


  buf

  (
    n1523_i2,
    g1399_n_spl_
  );


  buf

  (
    n464_i2,
    g1400_p_spl_
  );


  not

  (
    n1027_i2,
    g1401_n_spl_
  );


  not

  (
    n647_i2,
    g1402_n_spl_
  );


  not

  (
    n467_i2,
    g1403_n_spl_
  );


  buf

  (
    n2078_i2,
    g1407_p
  );


  not

  (
    n2079_i2,
    g1408_n
  );


  buf

  (
    n2178_i2,
    g1412_p
  );


  not

  (
    n2179_i2,
    g1413_n
  );


  buf

  (
    n2246_i2,
    g1417_p
  );


  not

  (
    n2247_i2,
    g1418_n
  );


  not

  (
    n2216_i2,
    g1422_p
  );


  not

  (
    n2217_i2,
    g1423_n
  );


  not

  (
    n2132_i2,
    g1427_p
  );


  not

  (
    n2133_i2,
    g1428_n
  );


  not

  (
    n2016_i2,
    g1432_p
  );


  not

  (
    n2017_i2,
    g1433_n
  );


  buf

  (
    n1946_i2,
    g1434_p
  );


  not

  (
    n1556_i2,
    g1438_n_spl_
  );


  not

  (
    n1752_i2,
    g1442_n_spl_
  );


  not

  (
    n1916_i2,
    g1446_n_spl_
  );


  not

  (
    n2048_i2,
    g1450_n_spl_
  );


  buf

  (
    n2102_i2,
    g1453_n_spl_
  );


  buf

  (
    n1226_i2,
    g1477_p_spl_
  );


  buf

  (
    n1986_i2,
    g1489_n_spl_
  );


  buf

  (
    n1838_i2,
    g1501_n_spl_
  );


  buf

  (
    n1658_i2,
    g1513_n_spl_
  );


  buf

  (
    n1123_i2,
    g1515_p_spl_
  );


  not

  (
    n1526_i2,
    g1519_n_spl_
  );


  not

  (
    n1722_i2,
    g1523_n_spl_
  );


  buf

  (
    n1808_i2,
    g1534_n_spl_
  );


  buf

  (
    n1628_i2,
    g1546_n_spl_
  );


  buf

  (
    n703_i2,
    g1577_p_spl_
  );


  buf

  (
    n483_i2,
    g1593_p_spl_
  );


  buf

  (
    n1583_i2,
    g1594_p
  );


  buf

  (
    n1787_i2,
    g1595_p
  );


  buf

  (
    n1959_i2,
    g1596_p
  );


  buf

  (
    n2099_i2,
    g1597_p
  );


  buf

  (
    n2033_i2,
    g1598_p
  );


  buf

  (
    n1877_i2,
    g1599_p
  );


  buf

  (
    n1689_i2,
    g1600_p
  );


  buf

  (
    n1355_i2,
    g1617_p
  );


  buf

  (
    n1469_i2,
    g1626_p
  );


  not

  (
    n1238_i2,
    g1627_n
  );


  not

  (
    n1227_i2,
    g1628_n
  );


  buf

  (
    n1124_i2,
    g1629_p
  );


  buf

  (
    n704_i2,
    g1630_p_spl_
  );


  buf

  (
    n484_i2,
    g1631_p_spl_
  );


  not

  (
    n1338_i2,
    g1633_p
  );


  not

  (
    n1449_i2,
    g1635_p
  );


  not

  (
    n1558_i2,
    g1637_p
  );


  not

  (
    n1754_i2,
    g1639_p
  );


  not

  (
    n1918_i2,
    g1641_p
  );


  not

  (
    n2050_i2,
    g1643_p
  );


  buf

  (
    n2104_i2,
    g1645_p
  );


  buf

  (
    n1988_i2,
    g1647_p
  );


  buf

  (
    n1840_i2,
    g1649_p
  );


  buf

  (
    n1660_i2,
    g1651_p
  );


  not

  (
    n708_i2,
    g1652_n
  );


  not

  (
    n768_i2,
    g1687_p
  );


  buf

  (
    lo102_buf_i2,
    n2782_lo_p
  );


  buf

  (
    n1631_i2,
    g1691_p
  );


  not

  (
    n1632_i2,
    g1692_n
  );


  buf

  (
    n1811_i2,
    g1696_p
  );


  not

  (
    n1812_i2,
    g1697_n
  );


  not

  (
    n1889_i2,
    g1700_p
  );


  not

  (
    n1890_i2,
    g1701_n
  );


  not

  (
    n1725_i2,
    g1705_p
  );


  not

  (
    n1726_i2,
    g1706_n
  );


  not

  (
    n917_i2,
    g1776_p
  );


  not

  (
    n918_i2,
    g1777_n
  );


  not

  (
    n1003_i2,
    g1814_p
  );


  not

  (
    n1004_i2,
    g1815_n
  );


  not

  (
    n1097_i2,
    g1851_p
  );


  not

  (
    n1098_i2,
    g1852_n
  );


  not

  (
    n1199_i2,
    g1880_p
  );


  not

  (
    n1200_i2,
    g1881_n
  );


  not

  (
    n1309_i2,
    g1901_p
  );


  not

  (
    n1310_i2,
    g1902_n
  );


  not

  (
    n1420_i2,
    g1914_p
  );


  not

  (
    n1421_i2,
    g1915_n
  );


  not

  (
    n1529_i2,
    g1919_p
  );


  not

  (
    n1530_i2,
    g1920_n
  );


  buf

  (
    n839_i2,
    g1924_n
  );


  buf

  (
    n840_i2,
    g1925_p
  );


  buf

  (
    n577_i2,
    g1975_n_spl_
  );


  buf

  (
    n623_i2,
    g1997_n_spl_
  );


  buf

  (
    n677_i2,
    g2019_n_spl_
  );


  buf

  (
    n739_i2,
    g2041_n_spl_
  );


  buf

  (
    n809_i2,
    g2063_n_spl_
  );


  buf

  (
    n887_i2,
    g2085_n_spl_
  );


  buf

  (
    n973_i2,
    g2107_n_spl_
  );


  buf

  (
    n1067_i2,
    g2129_n_spl_
  );


  buf

  (
    n1169_i2,
    g2151_n_spl_
  );


  buf

  (
    n1279_i2,
    g2173_n_spl_
  );


  buf

  (
    n1390_i2,
    g2189_n_spl_
  );


  buf

  (
    n1499_i2,
    g2200_n_spl_
  );


  buf

  (
    n539_i2,
    g2212_n_spl_
  );


  buf

  (
    lo082_buf_i2,
    G21_p_spl_11
  );


  buf

  (
    n555_i2,
    g2213_p
  );


  buf

  (
    n601_i2,
    g2214_p
  );


  buf

  (
    n655_i2,
    g2215_p
  );


  buf

  (
    n717_i2,
    g2216_p
  );


  buf

  (
    n787_i2,
    g2217_p
  );


  buf

  (
    n865_i2,
    g2218_p
  );


  buf

  (
    n951_i2,
    g2219_p
  );


  buf

  (
    n1045_i2,
    g2220_p
  );


  buf

  (
    n1147_i2,
    g2221_p
  );


  buf

  (
    n1257_i2,
    g2222_p
  );


  buf

  (
    n1374_i2,
    g2223_p
  );


  buf

  (
    n1488_i2,
    g2224_p
  );


  buf

  (
    n1602_i2,
    g2225_p
  );


  buf

  (
    n517_i2,
    g2226_p
  );


  buf

  (
    n1603_i2,
    g2227_p
  );


  not

  (
    n509_i2,
    g2231_p
  );


  not

  (
    n510_i2,
    g2232_n
  );


  buf

  (
    n579_i2,
    g2234_p
  );


  buf

  (
    n625_i2,
    g2236_p
  );


  buf

  (
    n679_i2,
    g2238_p
  );


  buf

  (
    n741_i2,
    g2240_p
  );


  buf

  (
    n811_i2,
    g2242_p
  );


  buf

  (
    n889_i2,
    g2244_p
  );


  buf

  (
    n975_i2,
    g2246_p
  );


  buf

  (
    n1069_i2,
    g2248_p
  );


  buf

  (
    n1171_i2,
    g2250_p
  );


  buf

  (
    n1281_i2,
    g2252_p
  );


  buf

  (
    n1392_i2,
    g2254_p
  );


  buf

  (
    n1501_i2,
    g2256_p
  );


  buf

  (
    n541_i2,
    g2258_p
  );


  buf

  (
    n1946_o2_p_spl_,
    n1946_o2_p
  );


  buf

  (
    n2016_o2_p_spl_,
    n2016_o2_p
  );


  buf

  (
    n2016_o2_n_spl_,
    n2016_o2_n
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g433_n_spl_,
    g433_n
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    n2078_o2_n_spl_,
    n2078_o2_n
  );


  buf

  (
    n2078_o2_p_spl_,
    n2078_o2_p
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g443_p_spl_,
    g443_p
  );


  buf

  (
    n2863_lo_p_spl_,
    n2863_lo_p
  );


  buf

  (
    n2863_lo_p_spl_0,
    n2863_lo_p_spl_
  );


  buf

  (
    n2863_lo_p_spl_00,
    n2863_lo_p_spl_0
  );


  buf

  (
    n2863_lo_p_spl_01,
    n2863_lo_p_spl_0
  );


  buf

  (
    n2863_lo_p_spl_1,
    n2863_lo_p_spl_
  );


  buf

  (
    n2863_lo_p_spl_10,
    n2863_lo_p_spl_1
  );


  buf

  (
    n2863_lo_n_spl_,
    n2863_lo_n
  );


  buf

  (
    n2863_lo_n_spl_0,
    n2863_lo_n_spl_
  );


  buf

  (
    n2863_lo_n_spl_00,
    n2863_lo_n_spl_0
  );


  buf

  (
    n2863_lo_n_spl_01,
    n2863_lo_n_spl_0
  );


  buf

  (
    n2863_lo_n_spl_1,
    n2863_lo_n_spl_
  );


  buf

  (
    n2863_lo_n_spl_10,
    n2863_lo_n_spl_1
  );


  buf

  (
    n2132_o2_p_spl_,
    n2132_o2_p
  );


  buf

  (
    n2132_o2_n_spl_,
    n2132_o2_n
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    n2178_o2_n_spl_,
    n2178_o2_n
  );


  buf

  (
    n2178_o2_p_spl_,
    n2178_o2_p
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g463_p_spl_,
    g463_p
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g463_n_spl_,
    g463_n
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g466_p_spl_,
    g466_p
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g466_n_spl_,
    g466_n
  );


  buf

  (
    g467_n_spl_,
    g467_n
  );


  buf

  (
    g467_p_spl_,
    g467_p
  );


  buf

  (
    g460_n_spl_,
    g460_n
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g470_n_spl_,
    g470_n
  );


  buf

  (
    g470_p_spl_,
    g470_p
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    n2635_lo_p_spl_,
    n2635_lo_p
  );


  buf

  (
    n2851_lo_p_spl_,
    n2851_lo_p
  );


  buf

  (
    n2851_lo_p_spl_0,
    n2851_lo_p_spl_
  );


  buf

  (
    n2851_lo_p_spl_1,
    n2851_lo_p_spl_
  );


  buf

  (
    n2635_lo_n_spl_,
    n2635_lo_n
  );


  buf

  (
    n2851_lo_n_spl_,
    n2851_lo_n
  );


  buf

  (
    n2851_lo_n_spl_0,
    n2851_lo_n_spl_
  );


  buf

  (
    n2851_lo_n_spl_1,
    n2851_lo_n_spl_
  );


  buf

  (
    n2216_o2_p_spl_,
    n2216_o2_p
  );


  buf

  (
    n2216_o2_n_spl_,
    n2216_o2_n
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g482_n_spl_,
    g482_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g487_p_spl_,
    g487_p
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g490_p_spl_,
    g490_p
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g490_n_spl_,
    g490_n
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g491_p_spl_,
    g491_p
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    n2647_lo_p_spl_,
    n2647_lo_p
  );


  buf

  (
    n2647_lo_n_spl_,
    n2647_lo_n
  );


  buf

  (
    n2246_o2_n_spl_,
    n2246_o2_n
  );


  buf

  (
    n2246_o2_p_spl_,
    n2246_o2_p
  );


  buf

  (
    g502_n_spl_,
    g502_n
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g502_p_spl_,
    g502_p
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g504_n_spl_,
    g504_n
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g501_n_spl_,
    g501_n
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g501_p_spl_,
    g501_p
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g507_n_spl_,
    g507_n
  );


  buf

  (
    g507_p_spl_,
    g507_p
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g510_n_spl_,
    g510_n
  );


  buf

  (
    g510_p_spl_,
    g510_p
  );


  buf

  (
    g499_n_spl_,
    g499_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g513_n_spl_,
    g513_n
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g498_n_spl_,
    g498_n
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g498_p_spl_,
    g498_p
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    g516_n_spl_,
    g516_n
  );


  buf

  (
    g516_p_spl_,
    g516_p
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g519_p_spl_,
    g519_p
  );


  buf

  (
    n2659_lo_p_spl_,
    n2659_lo_p
  );


  buf

  (
    n2659_lo_n_spl_,
    n2659_lo_n
  );


  buf

  (
    n2671_lo_p_spl_,
    n2671_lo_p
  );


  buf

  (
    n2671_lo_p_spl_0,
    n2671_lo_p_spl_
  );


  buf

  (
    n2671_lo_n_spl_,
    n2671_lo_n
  );


  buf

  (
    n2671_lo_n_spl_0,
    n2671_lo_n_spl_
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g528_p_spl_,
    g528_p
  );


  buf

  (
    g529_n_spl_,
    g529_n
  );


  buf

  (
    g529_p_spl_,
    g529_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    g526_p_spl_,
    g526_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g532_n_spl_,
    g532_n
  );


  buf

  (
    g532_p_spl_,
    g532_p
  );


  buf

  (
    g525_n_spl_,
    g525_n
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g525_p_spl_,
    g525_p
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g538_n_spl_,
    g538_n
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    g543_n_spl_,
    g543_n
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g549_n_spl_,
    g549_n
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g555_n_spl_,
    g555_n
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g548_n_spl_,
    g548_n
  );


  buf

  (
    g557_p_spl_,
    g557_p
  );


  buf

  (
    g548_p_spl_,
    g548_p
  );


  buf

  (
    g557_n_spl_,
    g557_n
  );


  buf

  (
    g558_n_spl_,
    g558_n
  );


  buf

  (
    g558_p_spl_,
    g558_p
  );


  buf

  (
    g547_p_spl_,
    g547_p
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g561_p_spl_,
    g561_p
  );


  buf

  (
    g564_n_spl_,
    g564_n
  );


  buf

  (
    g565_n_spl_,
    g565_n
  );


  buf

  (
    g564_p_spl_,
    g564_p
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g566_n_spl_,
    g566_n
  );


  buf

  (
    g570_n_spl_,
    g570_n
  );


  buf

  (
    n2848_lo_p_spl_,
    n2848_lo_p
  );


  buf

  (
    n2848_lo_p_spl_0,
    n2848_lo_p_spl_
  );


  buf

  (
    n2848_lo_p_spl_00,
    n2848_lo_p_spl_0
  );


  buf

  (
    n2848_lo_p_spl_000,
    n2848_lo_p_spl_00
  );


  buf

  (
    n2848_lo_p_spl_001,
    n2848_lo_p_spl_00
  );


  buf

  (
    n2848_lo_p_spl_01,
    n2848_lo_p_spl_0
  );


  buf

  (
    n2848_lo_p_spl_010,
    n2848_lo_p_spl_01
  );


  buf

  (
    n2848_lo_p_spl_011,
    n2848_lo_p_spl_01
  );


  buf

  (
    n2848_lo_p_spl_1,
    n2848_lo_p_spl_
  );


  buf

  (
    n2848_lo_p_spl_10,
    n2848_lo_p_spl_1
  );


  buf

  (
    n2848_lo_p_spl_11,
    n2848_lo_p_spl_1
  );


  buf

  (
    n4908_o2_p_spl_,
    n4908_o2_p
  );


  buf

  (
    n2848_lo_n_spl_,
    n2848_lo_n
  );


  buf

  (
    n2848_lo_n_spl_0,
    n2848_lo_n_spl_
  );


  buf

  (
    n2848_lo_n_spl_00,
    n2848_lo_n_spl_0
  );


  buf

  (
    n2848_lo_n_spl_000,
    n2848_lo_n_spl_00
  );


  buf

  (
    n2848_lo_n_spl_001,
    n2848_lo_n_spl_00
  );


  buf

  (
    n2848_lo_n_spl_01,
    n2848_lo_n_spl_0
  );


  buf

  (
    n2848_lo_n_spl_010,
    n2848_lo_n_spl_01
  );


  buf

  (
    n2848_lo_n_spl_011,
    n2848_lo_n_spl_01
  );


  buf

  (
    n2848_lo_n_spl_1,
    n2848_lo_n_spl_
  );


  buf

  (
    n2848_lo_n_spl_10,
    n2848_lo_n_spl_1
  );


  buf

  (
    n2848_lo_n_spl_11,
    n2848_lo_n_spl_1
  );


  buf

  (
    n4908_o2_n_spl_,
    n4908_o2_n
  );


  buf

  (
    n1124_o2_p_spl_,
    n1124_o2_p
  );


  buf

  (
    g575_n_spl_,
    g575_n
  );


  buf

  (
    g576_p_spl_,
    g576_p
  );


  buf

  (
    g575_p_spl_,
    g575_p
  );


  buf

  (
    g576_n_spl_,
    g576_n
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    n2860_lo_n_spl_,
    n2860_lo_n
  );


  buf

  (
    n2860_lo_n_spl_0,
    n2860_lo_n_spl_
  );


  buf

  (
    n2860_lo_n_spl_00,
    n2860_lo_n_spl_0
  );


  buf

  (
    n2860_lo_n_spl_000,
    n2860_lo_n_spl_00
  );


  buf

  (
    n2860_lo_n_spl_01,
    n2860_lo_n_spl_0
  );


  buf

  (
    n2860_lo_n_spl_1,
    n2860_lo_n_spl_
  );


  buf

  (
    n2860_lo_n_spl_10,
    n2860_lo_n_spl_1
  );


  buf

  (
    n2860_lo_n_spl_11,
    n2860_lo_n_spl_1
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    n4867_o2_p_spl_,
    n4867_o2_p
  );


  buf

  (
    n4867_o2_n_spl_,
    n4867_o2_n
  );


  buf

  (
    n1238_o2_n_spl_,
    n1238_o2_n
  );


  buf

  (
    n1338_o2_n_spl_,
    n1338_o2_n
  );


  buf

  (
    n1238_o2_p_spl_,
    n1238_o2_p
  );


  buf

  (
    n1338_o2_p_spl_,
    n1338_o2_p
  );


  buf

  (
    g584_n_spl_,
    g584_n
  );


  buf

  (
    g584_p_spl_,
    g584_p
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g583_p_spl_,
    g583_p
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g587_p_spl_,
    g587_p
  );


  buf

  (
    g582_n_spl_,
    g582_n
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g592_p_spl_,
    g592_p
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    n2860_lo_p_spl_,
    n2860_lo_p
  );


  buf

  (
    n2860_lo_p_spl_0,
    n2860_lo_p_spl_
  );


  buf

  (
    n2860_lo_p_spl_00,
    n2860_lo_p_spl_0
  );


  buf

  (
    n2860_lo_p_spl_01,
    n2860_lo_p_spl_0
  );


  buf

  (
    n2860_lo_p_spl_1,
    n2860_lo_p_spl_
  );


  buf

  (
    n2860_lo_p_spl_10,
    n2860_lo_p_spl_1
  );


  buf

  (
    n2860_lo_p_spl_11,
    n2860_lo_p_spl_1
  );


  buf

  (
    n4836_o2_p_spl_,
    n4836_o2_p
  );


  buf

  (
    n4836_o2_n_spl_,
    n4836_o2_n
  );


  buf

  (
    n1355_o2_n_spl_,
    n1355_o2_n
  );


  buf

  (
    n1449_o2_n_spl_,
    n1449_o2_n
  );


  buf

  (
    n1355_o2_p_spl_,
    n1355_o2_p
  );


  buf

  (
    n1449_o2_p_spl_,
    n1449_o2_p
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g604_p_spl_,
    g604_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g606_p_spl_,
    g606_p
  );


  buf

  (
    g607_n_spl_,
    g607_n
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g609_p_spl_,
    g609_p
  );


  buf

  (
    n4837_o2_p_spl_,
    n4837_o2_p
  );


  buf

  (
    n4837_o2_n_spl_,
    n4837_o2_n
  );


  buf

  (
    n1469_o2_n_spl_,
    n1469_o2_n
  );


  buf

  (
    n1558_o2_n_spl_,
    n1558_o2_n
  );


  buf

  (
    n1469_o2_p_spl_,
    n1469_o2_p
  );


  buf

  (
    n1558_o2_p_spl_,
    n1558_o2_p
  );


  buf

  (
    g615_n_spl_,
    g615_n
  );


  buf

  (
    g615_p_spl_,
    g615_p
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g618_n_spl_,
    g618_n
  );


  buf

  (
    g618_p_spl_,
    g618_p
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g620_n_spl_,
    g620_n
  );


  buf

  (
    g621_n_spl_,
    g621_n
  );


  buf

  (
    g621_p_spl_,
    g621_p
  );


  buf

  (
    g612_n_spl_,
    g612_n
  );


  buf

  (
    g623_p_spl_,
    g623_p
  );


  buf

  (
    g612_p_spl_,
    g612_p
  );


  buf

  (
    g623_n_spl_,
    g623_n
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g624_p_spl_,
    g624_p
  );


  buf

  (
    g611_n_spl_,
    g611_n
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    n6148_o2_p_spl_,
    n6148_o2_p
  );


  buf

  (
    n6148_o2_p_spl_0,
    n6148_o2_p_spl_
  );


  buf

  (
    n6148_o2_p_spl_00,
    n6148_o2_p_spl_0
  );


  buf

  (
    n6148_o2_p_spl_1,
    n6148_o2_p_spl_
  );


  buf

  (
    lo102_buf_o2_p_spl_,
    lo102_buf_o2_p
  );


  buf

  (
    lo102_buf_o2_p_spl_0,
    lo102_buf_o2_p_spl_
  );


  buf

  (
    lo102_buf_o2_p_spl_00,
    lo102_buf_o2_p_spl_0
  );


  buf

  (
    lo102_buf_o2_p_spl_000,
    lo102_buf_o2_p_spl_00
  );


  buf

  (
    lo102_buf_o2_p_spl_001,
    lo102_buf_o2_p_spl_00
  );


  buf

  (
    lo102_buf_o2_p_spl_01,
    lo102_buf_o2_p_spl_0
  );


  buf

  (
    lo102_buf_o2_p_spl_010,
    lo102_buf_o2_p_spl_01
  );


  buf

  (
    lo102_buf_o2_p_spl_011,
    lo102_buf_o2_p_spl_01
  );


  buf

  (
    lo102_buf_o2_p_spl_1,
    lo102_buf_o2_p_spl_
  );


  buf

  (
    lo102_buf_o2_p_spl_10,
    lo102_buf_o2_p_spl_1
  );


  buf

  (
    lo102_buf_o2_p_spl_100,
    lo102_buf_o2_p_spl_10
  );


  buf

  (
    lo102_buf_o2_p_spl_101,
    lo102_buf_o2_p_spl_10
  );


  buf

  (
    lo102_buf_o2_p_spl_11,
    lo102_buf_o2_p_spl_1
  );


  buf

  (
    lo102_buf_o2_p_spl_110,
    lo102_buf_o2_p_spl_11
  );


  buf

  (
    lo102_buf_o2_p_spl_111,
    lo102_buf_o2_p_spl_11
  );


  buf

  (
    n6148_o2_n_spl_,
    n6148_o2_n
  );


  buf

  (
    n6148_o2_n_spl_0,
    n6148_o2_n_spl_
  );


  buf

  (
    n6148_o2_n_spl_00,
    n6148_o2_n_spl_0
  );


  buf

  (
    n6148_o2_n_spl_1,
    n6148_o2_n_spl_
  );


  buf

  (
    lo102_buf_o2_n_spl_,
    lo102_buf_o2_n
  );


  buf

  (
    lo102_buf_o2_n_spl_0,
    lo102_buf_o2_n_spl_
  );


  buf

  (
    lo102_buf_o2_n_spl_00,
    lo102_buf_o2_n_spl_0
  );


  buf

  (
    lo102_buf_o2_n_spl_000,
    lo102_buf_o2_n_spl_00
  );


  buf

  (
    lo102_buf_o2_n_spl_001,
    lo102_buf_o2_n_spl_00
  );


  buf

  (
    lo102_buf_o2_n_spl_01,
    lo102_buf_o2_n_spl_0
  );


  buf

  (
    lo102_buf_o2_n_spl_010,
    lo102_buf_o2_n_spl_01
  );


  buf

  (
    lo102_buf_o2_n_spl_011,
    lo102_buf_o2_n_spl_01
  );


  buf

  (
    lo102_buf_o2_n_spl_1,
    lo102_buf_o2_n_spl_
  );


  buf

  (
    lo102_buf_o2_n_spl_10,
    lo102_buf_o2_n_spl_1
  );


  buf

  (
    lo102_buf_o2_n_spl_100,
    lo102_buf_o2_n_spl_10
  );


  buf

  (
    lo102_buf_o2_n_spl_101,
    lo102_buf_o2_n_spl_10
  );


  buf

  (
    lo102_buf_o2_n_spl_11,
    lo102_buf_o2_n_spl_1
  );


  buf

  (
    lo102_buf_o2_n_spl_110,
    lo102_buf_o2_n_spl_11
  );


  buf

  (
    lo102_buf_o2_n_spl_111,
    lo102_buf_o2_n_spl_11
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    n708_o2_n_spl_,
    n708_o2_n
  );


  buf

  (
    n768_o2_n_spl_,
    n768_o2_n
  );


  buf

  (
    n708_o2_p_spl_,
    n708_o2_p
  );


  buf

  (
    n768_o2_p_spl_,
    n768_o2_p
  );


  buf

  (
    g632_n_spl_,
    g632_n
  );


  buf

  (
    g632_p_spl_,
    g632_p
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g631_p_spl_,
    g631_p
  );


  buf

  (
    n4838_o2_p_spl_,
    n4838_o2_p
  );


  buf

  (
    n4838_o2_n_spl_,
    n4838_o2_n
  );


  buf

  (
    n1583_o2_n_spl_,
    n1583_o2_n
  );


  buf

  (
    n1660_o2_p_spl_,
    n1660_o2_p
  );


  buf

  (
    n1583_o2_p_spl_,
    n1583_o2_p
  );


  buf

  (
    n1660_o2_n_spl_,
    n1660_o2_n
  );


  buf

  (
    g642_n_spl_,
    g642_n
  );


  buf

  (
    g642_p_spl_,
    g642_p
  );


  buf

  (
    g641_n_spl_,
    g641_n
  );


  buf

  (
    g644_p_spl_,
    g644_p
  );


  buf

  (
    g641_p_spl_,
    g641_p
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g645_p_spl_,
    g645_p
  );


  buf

  (
    g640_n_spl_,
    g640_n
  );


  buf

  (
    g647_p_spl_,
    g647_p
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g639_n_spl_,
    g639_n
  );


  buf

  (
    g650_p_spl_,
    g650_p
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g650_n_spl_,
    g650_n
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g651_p_spl_,
    g651_p
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g637_n_spl_,
    g637_n
  );


  buf

  (
    g656_p_spl_,
    g656_p
  );


  buf

  (
    n2797_lo_p_spl_,
    n2797_lo_p
  );


  buf

  (
    n2797_lo_p_spl_0,
    n2797_lo_p_spl_
  );


  buf

  (
    n2797_lo_p_spl_00,
    n2797_lo_p_spl_0
  );


  buf

  (
    n2797_lo_p_spl_000,
    n2797_lo_p_spl_00
  );


  buf

  (
    n2797_lo_p_spl_001,
    n2797_lo_p_spl_00
  );


  buf

  (
    n2797_lo_p_spl_01,
    n2797_lo_p_spl_0
  );


  buf

  (
    n2797_lo_p_spl_010,
    n2797_lo_p_spl_01
  );


  buf

  (
    n2797_lo_p_spl_011,
    n2797_lo_p_spl_01
  );


  buf

  (
    n2797_lo_p_spl_1,
    n2797_lo_p_spl_
  );


  buf

  (
    n2797_lo_p_spl_10,
    n2797_lo_p_spl_1
  );


  buf

  (
    n2797_lo_p_spl_100,
    n2797_lo_p_spl_10
  );


  buf

  (
    n2797_lo_p_spl_101,
    n2797_lo_p_spl_10
  );


  buf

  (
    n2797_lo_p_spl_11,
    n2797_lo_p_spl_1
  );


  buf

  (
    n2797_lo_p_spl_110,
    n2797_lo_p_spl_11
  );


  buf

  (
    n2797_lo_p_spl_111,
    n2797_lo_p_spl_11
  );


  buf

  (
    n2797_lo_n_spl_,
    n2797_lo_n
  );


  buf

  (
    n2797_lo_n_spl_0,
    n2797_lo_n_spl_
  );


  buf

  (
    n2797_lo_n_spl_00,
    n2797_lo_n_spl_0
  );


  buf

  (
    n2797_lo_n_spl_000,
    n2797_lo_n_spl_00
  );


  buf

  (
    n2797_lo_n_spl_001,
    n2797_lo_n_spl_00
  );


  buf

  (
    n2797_lo_n_spl_01,
    n2797_lo_n_spl_0
  );


  buf

  (
    n2797_lo_n_spl_010,
    n2797_lo_n_spl_01
  );


  buf

  (
    n2797_lo_n_spl_011,
    n2797_lo_n_spl_01
  );


  buf

  (
    n2797_lo_n_spl_1,
    n2797_lo_n_spl_
  );


  buf

  (
    n2797_lo_n_spl_10,
    n2797_lo_n_spl_1
  );


  buf

  (
    n2797_lo_n_spl_100,
    n2797_lo_n_spl_10
  );


  buf

  (
    n2797_lo_n_spl_101,
    n2797_lo_n_spl_10
  );


  buf

  (
    n2797_lo_n_spl_11,
    n2797_lo_n_spl_1
  );


  buf

  (
    g636_n_spl_,
    g636_n
  );


  buf

  (
    g659_p_spl_,
    g659_p
  );


  buf

  (
    g635_p_spl_,
    g635_p
  );


  buf

  (
    n6053_o2_p_spl_,
    n6053_o2_p
  );


  buf

  (
    n6053_o2_p_spl_0,
    n6053_o2_p_spl_
  );


  buf

  (
    n6053_o2_p_spl_00,
    n6053_o2_p_spl_0
  );


  buf

  (
    n6053_o2_p_spl_1,
    n6053_o2_p_spl_
  );


  buf

  (
    n6053_o2_n_spl_,
    n6053_o2_n
  );


  buf

  (
    n6053_o2_n_spl_0,
    n6053_o2_n_spl_
  );


  buf

  (
    n6053_o2_n_spl_00,
    n6053_o2_n_spl_0
  );


  buf

  (
    n6053_o2_n_spl_1,
    n6053_o2_n_spl_
  );


  buf

  (
    n839_o2_p_spl_,
    n839_o2_p
  );


  buf

  (
    n839_o2_n_spl_,
    n839_o2_n
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    g664_p_spl_,
    g664_p
  );


  buf

  (
    g663_p_spl_,
    g663_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g665_n_spl_,
    g665_n
  );


  buf

  (
    g665_p_spl_,
    g665_p
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    g667_p_spl_,
    g667_p
  );


  buf

  (
    g662_p_spl_,
    g662_p
  );


  buf

  (
    g667_n_spl_,
    g667_n
  );


  buf

  (
    g668_n_spl_,
    g668_n
  );


  buf

  (
    g668_p_spl_,
    g668_p
  );


  buf

  (
    g670_p_spl_,
    g670_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    lo002_buf_o2_p_spl_,
    lo002_buf_o2_p
  );


  buf

  (
    lo002_buf_o2_p_spl_0,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    lo002_buf_o2_p_spl_00,
    lo002_buf_o2_p_spl_0
  );


  buf

  (
    lo002_buf_o2_p_spl_1,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    lo082_buf_o2_p_spl_,
    lo082_buf_o2_p
  );


  buf

  (
    lo082_buf_o2_p_spl_0,
    lo082_buf_o2_p_spl_
  );


  buf

  (
    lo002_buf_o2_n_spl_,
    lo002_buf_o2_n
  );


  buf

  (
    lo002_buf_o2_n_spl_0,
    lo002_buf_o2_n_spl_
  );


  buf

  (
    lo002_buf_o2_n_spl_00,
    lo002_buf_o2_n_spl_0
  );


  buf

  (
    lo002_buf_o2_n_spl_1,
    lo002_buf_o2_n_spl_
  );


  buf

  (
    lo082_buf_o2_n_spl_,
    lo082_buf_o2_n
  );


  buf

  (
    lo082_buf_o2_n_spl_0,
    lo082_buf_o2_n_spl_
  );


  buf

  (
    n509_o2_p_spl_,
    n509_o2_p
  );


  buf

  (
    n509_o2_n_spl_,
    n509_o2_n
  );


  buf

  (
    g661_p_spl_,
    g661_p
  );


  buf

  (
    n4839_o2_p_spl_,
    n4839_o2_p
  );


  buf

  (
    n4839_o2_n_spl_,
    n4839_o2_n
  );


  buf

  (
    n4840_o2_p_spl_,
    n4840_o2_p
  );


  buf

  (
    n4840_o2_p_spl_0,
    n4840_o2_p_spl_
  );


  buf

  (
    lo118_buf_o2_p_spl_,
    lo118_buf_o2_p
  );


  buf

  (
    lo118_buf_o2_p_spl_0,
    lo118_buf_o2_p_spl_
  );


  buf

  (
    lo118_buf_o2_p_spl_00,
    lo118_buf_o2_p_spl_0
  );


  buf

  (
    lo118_buf_o2_p_spl_000,
    lo118_buf_o2_p_spl_00
  );


  buf

  (
    lo118_buf_o2_p_spl_01,
    lo118_buf_o2_p_spl_0
  );


  buf

  (
    lo118_buf_o2_p_spl_1,
    lo118_buf_o2_p_spl_
  );


  buf

  (
    lo118_buf_o2_p_spl_10,
    lo118_buf_o2_p_spl_1
  );


  buf

  (
    lo118_buf_o2_p_spl_11,
    lo118_buf_o2_p_spl_1
  );


  buf

  (
    n4840_o2_n_spl_,
    n4840_o2_n
  );


  buf

  (
    n4840_o2_n_spl_0,
    n4840_o2_n_spl_
  );


  buf

  (
    lo118_buf_o2_n_spl_,
    lo118_buf_o2_n
  );


  buf

  (
    lo118_buf_o2_n_spl_0,
    lo118_buf_o2_n_spl_
  );


  buf

  (
    lo118_buf_o2_n_spl_00,
    lo118_buf_o2_n_spl_0
  );


  buf

  (
    lo118_buf_o2_n_spl_000,
    lo118_buf_o2_n_spl_00
  );


  buf

  (
    lo118_buf_o2_n_spl_01,
    lo118_buf_o2_n_spl_0
  );


  buf

  (
    lo118_buf_o2_n_spl_1,
    lo118_buf_o2_n_spl_
  );


  buf

  (
    lo118_buf_o2_n_spl_10,
    lo118_buf_o2_n_spl_1
  );


  buf

  (
    lo118_buf_o2_n_spl_11,
    lo118_buf_o2_n_spl_1
  );


  buf

  (
    n1689_o2_n_spl_,
    n1689_o2_n
  );


  buf

  (
    n1754_o2_n_spl_,
    n1754_o2_n
  );


  buf

  (
    n1689_o2_p_spl_,
    n1689_o2_p
  );


  buf

  (
    n1754_o2_p_spl_,
    n1754_o2_p
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g680_n_spl_,
    g680_n
  );


  buf

  (
    g683_p_spl_,
    g683_p
  );


  buf

  (
    g680_p_spl_,
    g680_p
  );


  buf

  (
    g683_n_spl_,
    g683_n
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g684_p_spl_,
    g684_p
  );


  buf

  (
    g679_n_spl_,
    g679_n
  );


  buf

  (
    g686_p_spl_,
    g686_p
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g686_n_spl_,
    g686_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g689_p_spl_,
    g689_p
  );


  buf

  (
    g678_p_spl_,
    g678_p
  );


  buf

  (
    g689_n_spl_,
    g689_n
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g677_n_spl_,
    g677_n
  );


  buf

  (
    g692_p_spl_,
    g692_p
  );


  buf

  (
    g677_p_spl_,
    g677_p
  );


  buf

  (
    g692_n_spl_,
    g692_n
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g695_p_spl_,
    g695_p
  );


  buf

  (
    g676_p_spl_,
    g676_p
  );


  buf

  (
    g695_n_spl_,
    g695_n
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    g698_p_spl_,
    g698_p
  );


  buf

  (
    g673_p_spl_,
    g673_p
  );


  buf

  (
    g672_p_spl_,
    g672_p
  );


  buf

  (
    n2809_lo_p_spl_,
    n2809_lo_p
  );


  buf

  (
    n2809_lo_p_spl_0,
    n2809_lo_p_spl_
  );


  buf

  (
    n2809_lo_p_spl_00,
    n2809_lo_p_spl_0
  );


  buf

  (
    n2809_lo_p_spl_000,
    n2809_lo_p_spl_00
  );


  buf

  (
    n2809_lo_p_spl_001,
    n2809_lo_p_spl_00
  );


  buf

  (
    n2809_lo_p_spl_01,
    n2809_lo_p_spl_0
  );


  buf

  (
    n2809_lo_p_spl_010,
    n2809_lo_p_spl_01
  );


  buf

  (
    n2809_lo_p_spl_011,
    n2809_lo_p_spl_01
  );


  buf

  (
    n2809_lo_p_spl_1,
    n2809_lo_p_spl_
  );


  buf

  (
    n2809_lo_p_spl_10,
    n2809_lo_p_spl_1
  );


  buf

  (
    n2809_lo_p_spl_100,
    n2809_lo_p_spl_10
  );


  buf

  (
    n2809_lo_p_spl_11,
    n2809_lo_p_spl_1
  );


  buf

  (
    n2809_lo_n_spl_,
    n2809_lo_n
  );


  buf

  (
    n2809_lo_n_spl_0,
    n2809_lo_n_spl_
  );


  buf

  (
    n2809_lo_n_spl_00,
    n2809_lo_n_spl_0
  );


  buf

  (
    n2809_lo_n_spl_000,
    n2809_lo_n_spl_00
  );


  buf

  (
    n2809_lo_n_spl_001,
    n2809_lo_n_spl_00
  );


  buf

  (
    n2809_lo_n_spl_01,
    n2809_lo_n_spl_0
  );


  buf

  (
    n2809_lo_n_spl_010,
    n2809_lo_n_spl_01
  );


  buf

  (
    n2809_lo_n_spl_1,
    n2809_lo_n_spl_
  );


  buf

  (
    n2809_lo_n_spl_10,
    n2809_lo_n_spl_1
  );


  buf

  (
    n2809_lo_n_spl_11,
    n2809_lo_n_spl_1
  );


  buf

  (
    n2734_lo_p_spl_,
    n2734_lo_p
  );


  buf

  (
    n2734_lo_p_spl_0,
    n2734_lo_p_spl_
  );


  buf

  (
    n2734_lo_p_spl_00,
    n2734_lo_p_spl_0
  );


  buf

  (
    n2734_lo_p_spl_000,
    n2734_lo_p_spl_00
  );


  buf

  (
    n2734_lo_p_spl_001,
    n2734_lo_p_spl_00
  );


  buf

  (
    n2734_lo_p_spl_01,
    n2734_lo_p_spl_0
  );


  buf

  (
    n2734_lo_p_spl_010,
    n2734_lo_p_spl_01
  );


  buf

  (
    n2734_lo_p_spl_011,
    n2734_lo_p_spl_01
  );


  buf

  (
    n2734_lo_p_spl_1,
    n2734_lo_p_spl_
  );


  buf

  (
    n2734_lo_p_spl_10,
    n2734_lo_p_spl_1
  );


  buf

  (
    n2734_lo_p_spl_100,
    n2734_lo_p_spl_10
  );


  buf

  (
    n2734_lo_p_spl_101,
    n2734_lo_p_spl_10
  );


  buf

  (
    n2734_lo_p_spl_11,
    n2734_lo_p_spl_1
  );


  buf

  (
    n2734_lo_p_spl_110,
    n2734_lo_p_spl_11
  );


  buf

  (
    n2734_lo_p_spl_111,
    n2734_lo_p_spl_11
  );


  buf

  (
    n2734_lo_n_spl_,
    n2734_lo_n
  );


  buf

  (
    n2734_lo_n_spl_0,
    n2734_lo_n_spl_
  );


  buf

  (
    n2734_lo_n_spl_00,
    n2734_lo_n_spl_0
  );


  buf

  (
    n2734_lo_n_spl_000,
    n2734_lo_n_spl_00
  );


  buf

  (
    n2734_lo_n_spl_001,
    n2734_lo_n_spl_00
  );


  buf

  (
    n2734_lo_n_spl_01,
    n2734_lo_n_spl_0
  );


  buf

  (
    n2734_lo_n_spl_010,
    n2734_lo_n_spl_01
  );


  buf

  (
    n2734_lo_n_spl_011,
    n2734_lo_n_spl_01
  );


  buf

  (
    n2734_lo_n_spl_1,
    n2734_lo_n_spl_
  );


  buf

  (
    n2734_lo_n_spl_10,
    n2734_lo_n_spl_1
  );


  buf

  (
    n2734_lo_n_spl_100,
    n2734_lo_n_spl_10
  );


  buf

  (
    n2734_lo_n_spl_101,
    n2734_lo_n_spl_10
  );


  buf

  (
    n2734_lo_n_spl_11,
    n2734_lo_n_spl_1
  );


  buf

  (
    n2734_lo_n_spl_110,
    n2734_lo_n_spl_11
  );


  buf

  (
    n2734_lo_n_spl_111,
    n2734_lo_n_spl_11
  );


  buf

  (
    n2099_o2_n_spl_,
    n2099_o2_n
  );


  buf

  (
    n2104_o2_p_spl_,
    n2104_o2_p
  );


  buf

  (
    n2099_o2_p_spl_,
    n2099_o2_p
  );


  buf

  (
    n2104_o2_n_spl_,
    n2104_o2_n
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    n4847_o2_p_spl_,
    n4847_o2_p
  );


  buf

  (
    n4847_o2_p_spl_0,
    n4847_o2_p_spl_
  );


  buf

  (
    n4847_o2_p_spl_1,
    n4847_o2_p_spl_
  );


  buf

  (
    lo110_buf_o2_p_spl_,
    lo110_buf_o2_p
  );


  buf

  (
    lo110_buf_o2_p_spl_0,
    lo110_buf_o2_p_spl_
  );


  buf

  (
    lo110_buf_o2_p_spl_1,
    lo110_buf_o2_p_spl_
  );


  buf

  (
    n4847_o2_n_spl_,
    n4847_o2_n
  );


  buf

  (
    n4847_o2_n_spl_0,
    n4847_o2_n_spl_
  );


  buf

  (
    lo110_buf_o2_n_spl_,
    lo110_buf_o2_n
  );


  buf

  (
    lo110_buf_o2_n_spl_0,
    lo110_buf_o2_n_spl_
  );


  buf

  (
    lo110_buf_o2_n_spl_1,
    lo110_buf_o2_n_spl_
  );


  buf

  (
    g709_n_spl_,
    g709_n
  );


  buf

  (
    g709_p_spl_,
    g709_p
  );


  buf

  (
    g710_n_spl_,
    g710_n
  );


  buf

  (
    g712_p_spl_,
    g712_p
  );


  buf

  (
    g710_p_spl_,
    g710_p
  );


  buf

  (
    g712_n_spl_,
    g712_n
  );


  buf

  (
    g713_n_spl_,
    g713_n
  );


  buf

  (
    g713_p_spl_,
    g713_p
  );


  buf

  (
    n4848_o2_p_spl_,
    n4848_o2_p
  );


  buf

  (
    n4848_o2_p_spl_0,
    n4848_o2_p_spl_
  );


  buf

  (
    n4848_o2_n_spl_,
    n4848_o2_n
  );


  buf

  (
    n4848_o2_n_spl_0,
    n4848_o2_n_spl_
  );


  buf

  (
    n4849_o2_p_spl_,
    n4849_o2_p
  );


  buf

  (
    n4849_o2_p_spl_0,
    n4849_o2_p_spl_
  );


  buf

  (
    n4849_o2_p_spl_1,
    n4849_o2_p_spl_
  );


  buf

  (
    n4849_o2_n_spl_,
    n4849_o2_n
  );


  buf

  (
    n4849_o2_n_spl_0,
    n4849_o2_n_spl_
  );


  buf

  (
    g716_n_spl_,
    g716_n
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g716_p_spl_,
    g716_p
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


  buf

  (
    g718_p_spl_,
    g718_p
  );


  buf

  (
    g715_n_spl_,
    g715_n
  );


  buf

  (
    g720_p_spl_,
    g720_p
  );


  buf

  (
    g715_p_spl_,
    g715_p
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g721_n_spl_,
    g721_n
  );


  buf

  (
    g721_p_spl_,
    g721_p
  );


  buf

  (
    g714_n_spl_,
    g714_n
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    lo114_buf_o2_p_spl_,
    lo114_buf_o2_p
  );


  buf

  (
    lo114_buf_o2_p_spl_0,
    lo114_buf_o2_p_spl_
  );


  buf

  (
    lo114_buf_o2_p_spl_00,
    lo114_buf_o2_p_spl_0
  );


  buf

  (
    lo114_buf_o2_p_spl_01,
    lo114_buf_o2_p_spl_0
  );


  buf

  (
    lo114_buf_o2_p_spl_1,
    lo114_buf_o2_p_spl_
  );


  buf

  (
    lo114_buf_o2_p_spl_10,
    lo114_buf_o2_p_spl_1
  );


  buf

  (
    lo114_buf_o2_n_spl_,
    lo114_buf_o2_n
  );


  buf

  (
    lo114_buf_o2_n_spl_0,
    lo114_buf_o2_n_spl_
  );


  buf

  (
    lo114_buf_o2_n_spl_00,
    lo114_buf_o2_n_spl_0
  );


  buf

  (
    lo114_buf_o2_n_spl_01,
    lo114_buf_o2_n_spl_0
  );


  buf

  (
    lo114_buf_o2_n_spl_1,
    lo114_buf_o2_n_spl_
  );


  buf

  (
    lo114_buf_o2_n_spl_10,
    lo114_buf_o2_n_spl_1
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g725_n_spl_,
    g725_n
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    g725_p_spl_,
    g725_p
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g728_n_spl_,
    g728_n
  );


  buf

  (
    g728_p_spl_,
    g728_p
  );


  buf

  (
    g731_n_spl_,
    g731_n
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g733_n_spl_,
    g733_n
  );


  buf

  (
    g733_p_spl_,
    g733_p
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g736_n_spl_,
    g736_n
  );


  buf

  (
    g736_p_spl_,
    g736_p
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    n1959_o2_n_spl_,
    n1959_o2_n
  );


  buf

  (
    n1988_o2_p_spl_,
    n1988_o2_p
  );


  buf

  (
    n1959_o2_p_spl_,
    n1959_o2_p
  );


  buf

  (
    n1988_o2_n_spl_,
    n1988_o2_n
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    g741_p_spl_,
    g741_p
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g743_n_spl_,
    g743_n
  );


  buf

  (
    n4844_o2_p_spl_,
    n4844_o2_p
  );


  buf

  (
    n4844_o2_p_spl_0,
    n4844_o2_p_spl_
  );


  buf

  (
    n4844_o2_p_spl_1,
    n4844_o2_p_spl_
  );


  buf

  (
    n4844_o2_n_spl_,
    n4844_o2_n
  );


  buf

  (
    n4844_o2_n_spl_0,
    n4844_o2_n_spl_
  );


  buf

  (
    g744_n_spl_,
    g744_n
  );


  buf

  (
    g744_p_spl_,
    g744_p
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g745_p_spl_,
    g745_p
  );


  buf

  (
    g747_n_spl_,
    g747_n
  );


  buf

  (
    g748_n_spl_,
    g748_n
  );


  buf

  (
    g748_p_spl_,
    g748_p
  );


  buf

  (
    n4845_o2_p_spl_,
    n4845_o2_p
  );


  buf

  (
    n4845_o2_p_spl_0,
    n4845_o2_p_spl_
  );


  buf

  (
    n4845_o2_n_spl_,
    n4845_o2_n
  );


  buf

  (
    n4845_o2_n_spl_0,
    n4845_o2_n_spl_
  );


  buf

  (
    n4846_o2_p_spl_,
    n4846_o2_p
  );


  buf

  (
    n4846_o2_p_spl_0,
    n4846_o2_p_spl_
  );


  buf

  (
    n4846_o2_p_spl_1,
    n4846_o2_p_spl_
  );


  buf

  (
    n4846_o2_n_spl_,
    n4846_o2_n
  );


  buf

  (
    n4846_o2_n_spl_0,
    n4846_o2_n_spl_
  );


  buf

  (
    n2033_o2_n_spl_,
    n2033_o2_n
  );


  buf

  (
    n2050_o2_n_spl_,
    n2050_o2_n
  );


  buf

  (
    n2033_o2_p_spl_,
    n2033_o2_p
  );


  buf

  (
    n2050_o2_p_spl_,
    n2050_o2_p
  );


  buf

  (
    g753_n_spl_,
    g753_n
  );


  buf

  (
    g753_p_spl_,
    g753_p
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g752_p_spl_,
    g752_p
  );


  buf

  (
    g755_n_spl_,
    g755_n
  );


  buf

  (
    g756_n_spl_,
    g756_n
  );


  buf

  (
    g756_p_spl_,
    g756_p
  );


  buf

  (
    g751_n_spl_,
    g751_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g751_p_spl_,
    g751_p
  );


  buf

  (
    g758_n_spl_,
    g758_n
  );


  buf

  (
    g759_n_spl_,
    g759_n
  );


  buf

  (
    g759_p_spl_,
    g759_p
  );


  buf

  (
    g750_n_spl_,
    g750_n
  );


  buf

  (
    g761_p_spl_,
    g761_p
  );


  buf

  (
    g750_p_spl_,
    g750_p
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g762_n_spl_,
    g762_n
  );


  buf

  (
    g762_p_spl_,
    g762_p
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    g764_p_spl_,
    g764_p
  );


  buf

  (
    g749_p_spl_,
    g749_p
  );


  buf

  (
    g764_n_spl_,
    g764_n
  );


  buf

  (
    g765_n_spl_,
    g765_n
  );


  buf

  (
    g765_p_spl_,
    g765_p
  );


  buf

  (
    g766_n_spl_,
    g766_n
  );


  buf

  (
    g768_p_spl_,
    g768_p
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g768_n_spl_,
    g768_n
  );


  buf

  (
    g769_n_spl_,
    g769_n
  );


  buf

  (
    g769_p_spl_,
    g769_p
  );


  buf

  (
    g774_n_spl_,
    g774_n
  );


  buf

  (
    g776_p_spl_,
    g776_p
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g776_n_spl_,
    g776_n
  );


  buf

  (
    g777_n_spl_,
    g777_n
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    g773_n_spl_,
    g773_n
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g773_p_spl_,
    g773_p
  );


  buf

  (
    g779_n_spl_,
    g779_n
  );


  buf

  (
    g780_n_spl_,
    g780_n
  );


  buf

  (
    g780_p_spl_,
    g780_p
  );


  buf

  (
    g772_n_spl_,
    g772_n
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    g772_p_spl_,
    g772_p
  );


  buf

  (
    g782_n_spl_,
    g782_n
  );


  buf

  (
    g783_n_spl_,
    g783_n
  );


  buf

  (
    g783_p_spl_,
    g783_p
  );


  buf

  (
    g771_n_spl_,
    g771_n
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    g771_p_spl_,
    g771_p
  );


  buf

  (
    g785_n_spl_,
    g785_n
  );


  buf

  (
    g786_n_spl_,
    g786_n
  );


  buf

  (
    g786_p_spl_,
    g786_p
  );


  buf

  (
    g770_n_spl_,
    g770_n
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g770_p_spl_,
    g770_p
  );


  buf

  (
    g788_n_spl_,
    g788_n
  );


  buf

  (
    n1787_o2_n_spl_,
    n1787_o2_n
  );


  buf

  (
    n1840_o2_p_spl_,
    n1840_o2_p
  );


  buf

  (
    n1787_o2_p_spl_,
    n1787_o2_p
  );


  buf

  (
    n1840_o2_n_spl_,
    n1840_o2_n
  );


  buf

  (
    g791_n_spl_,
    g791_n
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    g790_n_spl_,
    g790_n
  );


  buf

  (
    g793_p_spl_,
    g793_p
  );


  buf

  (
    g790_p_spl_,
    g790_p
  );


  buf

  (
    g793_n_spl_,
    g793_n
  );


  buf

  (
    n4841_o2_p_spl_,
    n4841_o2_p
  );


  buf

  (
    n4841_o2_p_spl_0,
    n4841_o2_p_spl_
  );


  buf

  (
    n4841_o2_n_spl_,
    n4841_o2_n
  );


  buf

  (
    n4841_o2_n_spl_0,
    n4841_o2_n_spl_
  );


  buf

  (
    g794_n_spl_,
    g794_n
  );


  buf

  (
    g794_p_spl_,
    g794_p
  );


  buf

  (
    g795_n_spl_,
    g795_n
  );


  buf

  (
    g797_p_spl_,
    g797_p
  );


  buf

  (
    g795_p_spl_,
    g795_p
  );


  buf

  (
    g797_n_spl_,
    g797_n
  );


  buf

  (
    g798_n_spl_,
    g798_n
  );


  buf

  (
    g798_p_spl_,
    g798_p
  );


  buf

  (
    n4842_o2_p_spl_,
    n4842_o2_p
  );


  buf

  (
    n4842_o2_n_spl_,
    n4842_o2_n
  );


  buf

  (
    n4842_o2_n_spl_0,
    n4842_o2_n_spl_
  );


  buf

  (
    n4843_o2_p_spl_,
    n4843_o2_p
  );


  buf

  (
    n4843_o2_p_spl_0,
    n4843_o2_p_spl_
  );


  buf

  (
    n4843_o2_p_spl_1,
    n4843_o2_p_spl_
  );


  buf

  (
    n4843_o2_n_spl_,
    n4843_o2_n
  );


  buf

  (
    n4843_o2_n_spl_0,
    n4843_o2_n_spl_
  );


  buf

  (
    n1877_o2_n_spl_,
    n1877_o2_n
  );


  buf

  (
    n1918_o2_n_spl_,
    n1918_o2_n
  );


  buf

  (
    n1877_o2_p_spl_,
    n1877_o2_p
  );


  buf

  (
    n1918_o2_p_spl_,
    n1918_o2_p
  );


  buf

  (
    g803_n_spl_,
    g803_n
  );


  buf

  (
    g803_p_spl_,
    g803_p
  );


  buf

  (
    g802_n_spl_,
    g802_n
  );


  buf

  (
    g805_p_spl_,
    g805_p
  );


  buf

  (
    g802_p_spl_,
    g802_p
  );


  buf

  (
    g805_n_spl_,
    g805_n
  );


  buf

  (
    g806_n_spl_,
    g806_n
  );


  buf

  (
    g806_p_spl_,
    g806_p
  );


  buf

  (
    g801_n_spl_,
    g801_n
  );


  buf

  (
    g808_p_spl_,
    g808_p
  );


  buf

  (
    g801_p_spl_,
    g801_p
  );


  buf

  (
    g808_n_spl_,
    g808_n
  );


  buf

  (
    g809_n_spl_,
    g809_n
  );


  buf

  (
    g809_p_spl_,
    g809_p
  );


  buf

  (
    g800_n_spl_,
    g800_n
  );


  buf

  (
    g811_p_spl_,
    g811_p
  );


  buf

  (
    g800_p_spl_,
    g800_p
  );


  buf

  (
    g811_n_spl_,
    g811_n
  );


  buf

  (
    g812_n_spl_,
    g812_n
  );


  buf

  (
    g812_p_spl_,
    g812_p
  );


  buf

  (
    g799_n_spl_,
    g799_n
  );


  buf

  (
    g814_p_spl_,
    g814_p
  );


  buf

  (
    g799_p_spl_,
    g799_p
  );


  buf

  (
    g814_n_spl_,
    g814_n
  );


  buf

  (
    g815_n_spl_,
    g815_n
  );


  buf

  (
    g815_p_spl_,
    g815_p
  );


  buf

  (
    g816_n_spl_,
    g816_n
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g816_p_spl_,
    g816_p
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g819_n_spl_,
    g819_n
  );


  buf

  (
    g819_p_spl_,
    g819_p
  );


  buf

  (
    g824_n_spl_,
    g824_n
  );


  buf

  (
    g826_p_spl_,
    g826_p
  );


  buf

  (
    g824_p_spl_,
    g824_p
  );


  buf

  (
    g826_n_spl_,
    g826_n
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g823_n_spl_,
    g823_n
  );


  buf

  (
    g829_p_spl_,
    g829_p
  );


  buf

  (
    g823_p_spl_,
    g823_p
  );


  buf

  (
    g829_n_spl_,
    g829_n
  );


  buf

  (
    g830_n_spl_,
    g830_n
  );


  buf

  (
    g830_p_spl_,
    g830_p
  );


  buf

  (
    g822_n_spl_,
    g822_n
  );


  buf

  (
    g832_p_spl_,
    g832_p
  );


  buf

  (
    g822_p_spl_,
    g822_p
  );


  buf

  (
    g832_n_spl_,
    g832_n
  );


  buf

  (
    g833_n_spl_,
    g833_n
  );


  buf

  (
    g833_p_spl_,
    g833_p
  );


  buf

  (
    g821_n_spl_,
    g821_n
  );


  buf

  (
    g835_p_spl_,
    g835_p
  );


  buf

  (
    g821_p_spl_,
    g821_p
  );


  buf

  (
    g835_n_spl_,
    g835_n
  );


  buf

  (
    g836_n_spl_,
    g836_n
  );


  buf

  (
    g836_p_spl_,
    g836_p
  );


  buf

  (
    g820_n_spl_,
    g820_n
  );


  buf

  (
    g838_p_spl_,
    g838_p
  );


  buf

  (
    g820_p_spl_,
    g820_p
  );


  buf

  (
    g838_n_spl_,
    g838_n
  );


  buf

  (
    g674_n_spl_,
    g674_n
  );


  buf

  (
    g701_p_spl_,
    g701_p
  );


  buf

  (
    g671_p_spl_,
    g671_p
  );


  buf

  (
    n6024_o2_p_spl_,
    n6024_o2_p
  );


  buf

  (
    n6024_o2_p_spl_0,
    n6024_o2_p_spl_
  );


  buf

  (
    n6024_o2_p_spl_00,
    n6024_o2_p_spl_0
  );


  buf

  (
    n6024_o2_p_spl_01,
    n6024_o2_p_spl_0
  );


  buf

  (
    n6024_o2_p_spl_1,
    n6024_o2_p_spl_
  );


  buf

  (
    n6024_o2_n_spl_,
    n6024_o2_n
  );


  buf

  (
    n6024_o2_n_spl_0,
    n6024_o2_n_spl_
  );


  buf

  (
    n6024_o2_n_spl_00,
    n6024_o2_n_spl_0
  );


  buf

  (
    n6024_o2_n_spl_1,
    n6024_o2_n_spl_
  );


  buf

  (
    n917_o2_p_spl_,
    n917_o2_p
  );


  buf

  (
    n917_o2_n_spl_,
    n917_o2_n
  );


  buf

  (
    g844_n_spl_,
    g844_n
  );


  buf

  (
    g845_p_spl_,
    g845_p
  );


  buf

  (
    g844_p_spl_,
    g844_p
  );


  buf

  (
    g845_n_spl_,
    g845_n
  );


  buf

  (
    g846_n_spl_,
    g846_n
  );


  buf

  (
    g846_p_spl_,
    g846_p
  );


  buf

  (
    g843_n_spl_,
    g843_n
  );


  buf

  (
    g848_p_spl_,
    g848_p
  );


  buf

  (
    g843_p_spl_,
    g843_p
  );


  buf

  (
    g848_n_spl_,
    g848_n
  );


  buf

  (
    g849_n_spl_,
    g849_n
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g842_n_spl_,
    g842_n
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g842_p_spl_,
    g842_p
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g852_n_spl_,
    g852_n
  );


  buf

  (
    g852_p_spl_,
    g852_p
  );


  buf

  (
    g841_n_spl_,
    g841_n
  );


  buf

  (
    g854_p_spl_,
    g854_p
  );


  buf

  (
    g841_p_spl_,
    g841_p
  );


  buf

  (
    g854_n_spl_,
    g854_n
  );


  buf

  (
    g855_n_spl_,
    g855_n
  );


  buf

  (
    g855_p_spl_,
    g855_p
  );


  buf

  (
    g702_p_spl_,
    g702_p
  );


  buf

  (
    n517_o2_n_spl_,
    n517_o2_n
  );


  buf

  (
    n541_o2_p_spl_,
    n541_o2_p
  );


  buf

  (
    n517_o2_p_spl_,
    n517_o2_p
  );


  buf

  (
    n541_o2_n_spl_,
    n541_o2_n
  );


  buf

  (
    g859_n_spl_,
    g859_n
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g858_n_spl_,
    g858_n
  );


  buf

  (
    g861_p_spl_,
    g861_p
  );


  buf

  (
    g858_p_spl_,
    g858_p
  );


  buf

  (
    g861_n_spl_,
    g861_n
  );


  buf

  (
    g862_n_spl_,
    g862_n
  );


  buf

  (
    g862_p_spl_,
    g862_p
  );


  buf

  (
    g857_p_spl_,
    g857_p
  );


  buf

  (
    g703_p_spl_,
    g703_p
  );


  buf

  (
    g864_p_spl_,
    g864_p
  );


  buf

  (
    g704_p_spl_,
    g704_p
  );


  buf

  (
    g840_p_spl_,
    g840_p
  );


  buf

  (
    g872_n_spl_,
    g872_n
  );


  buf

  (
    g874_p_spl_,
    g874_p
  );


  buf

  (
    g872_p_spl_,
    g872_p
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g875_p_spl_,
    g875_p
  );


  buf

  (
    g871_n_spl_,
    g871_n
  );


  buf

  (
    g877_p_spl_,
    g877_p
  );


  buf

  (
    g871_p_spl_,
    g871_p
  );


  buf

  (
    g877_n_spl_,
    g877_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g878_p_spl_,
    g878_p
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    g880_p_spl_,
    g880_p
  );


  buf

  (
    g870_p_spl_,
    g870_p
  );


  buf

  (
    g880_n_spl_,
    g880_n
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g883_p_spl_,
    g883_p
  );


  buf

  (
    g869_p_spl_,
    g869_p
  );


  buf

  (
    g883_n_spl_,
    g883_n
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g884_p_spl_,
    g884_p
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    n2746_lo_p_spl_,
    n2746_lo_p
  );


  buf

  (
    n2746_lo_p_spl_0,
    n2746_lo_p_spl_
  );


  buf

  (
    n2746_lo_p_spl_00,
    n2746_lo_p_spl_0
  );


  buf

  (
    n2746_lo_p_spl_000,
    n2746_lo_p_spl_00
  );


  buf

  (
    n2746_lo_p_spl_001,
    n2746_lo_p_spl_00
  );


  buf

  (
    n2746_lo_p_spl_01,
    n2746_lo_p_spl_0
  );


  buf

  (
    n2746_lo_p_spl_010,
    n2746_lo_p_spl_01
  );


  buf

  (
    n2746_lo_p_spl_011,
    n2746_lo_p_spl_01
  );


  buf

  (
    n2746_lo_p_spl_1,
    n2746_lo_p_spl_
  );


  buf

  (
    n2746_lo_p_spl_10,
    n2746_lo_p_spl_1
  );


  buf

  (
    n2746_lo_p_spl_100,
    n2746_lo_p_spl_10
  );


  buf

  (
    n2746_lo_p_spl_101,
    n2746_lo_p_spl_10
  );


  buf

  (
    n2746_lo_p_spl_11,
    n2746_lo_p_spl_1
  );


  buf

  (
    n2746_lo_p_spl_110,
    n2746_lo_p_spl_11
  );


  buf

  (
    n2746_lo_n_spl_,
    n2746_lo_n
  );


  buf

  (
    n2746_lo_n_spl_0,
    n2746_lo_n_spl_
  );


  buf

  (
    n2746_lo_n_spl_00,
    n2746_lo_n_spl_0
  );


  buf

  (
    n2746_lo_n_spl_000,
    n2746_lo_n_spl_00
  );


  buf

  (
    n2746_lo_n_spl_001,
    n2746_lo_n_spl_00
  );


  buf

  (
    n2746_lo_n_spl_01,
    n2746_lo_n_spl_0
  );


  buf

  (
    n2746_lo_n_spl_010,
    n2746_lo_n_spl_01
  );


  buf

  (
    n2746_lo_n_spl_011,
    n2746_lo_n_spl_01
  );


  buf

  (
    n2746_lo_n_spl_1,
    n2746_lo_n_spl_
  );


  buf

  (
    n2746_lo_n_spl_10,
    n2746_lo_n_spl_1
  );


  buf

  (
    n2746_lo_n_spl_100,
    n2746_lo_n_spl_10
  );


  buf

  (
    n2746_lo_n_spl_101,
    n2746_lo_n_spl_10
  );


  buf

  (
    n2746_lo_n_spl_11,
    n2746_lo_n_spl_1
  );


  buf

  (
    n2746_lo_n_spl_110,
    n2746_lo_n_spl_11
  );


  buf

  (
    n2746_lo_n_spl_111,
    n2746_lo_n_spl_11
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    lo006_buf_o2_p_spl_,
    lo006_buf_o2_p
  );


  buf

  (
    lo006_buf_o2_p_spl_0,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    lo006_buf_o2_p_spl_00,
    lo006_buf_o2_p_spl_0
  );


  buf

  (
    lo006_buf_o2_p_spl_1,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    lo006_buf_o2_n_spl_,
    lo006_buf_o2_n
  );


  buf

  (
    lo006_buf_o2_n_spl_0,
    lo006_buf_o2_n_spl_
  );


  buf

  (
    lo006_buf_o2_n_spl_1,
    lo006_buf_o2_n_spl_
  );


  buf

  (
    n555_o2_n_spl_,
    n555_o2_n
  );


  buf

  (
    n579_o2_p_spl_,
    n579_o2_p
  );


  buf

  (
    n555_o2_p_spl_,
    n555_o2_p
  );


  buf

  (
    n579_o2_n_spl_,
    n579_o2_n
  );


  buf

  (
    g894_n_spl_,
    g894_n
  );


  buf

  (
    g894_p_spl_,
    g894_p
  );


  buf

  (
    g893_n_spl_,
    g893_n
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g893_p_spl_,
    g893_p
  );


  buf

  (
    g896_n_spl_,
    g896_n
  );


  buf

  (
    g897_n_spl_,
    g897_n
  );


  buf

  (
    g897_p_spl_,
    g897_p
  );


  buf

  (
    g892_n_spl_,
    g892_n
  );


  buf

  (
    g899_p_spl_,
    g899_p
  );


  buf

  (
    g892_p_spl_,
    g892_p
  );


  buf

  (
    g899_n_spl_,
    g899_n
  );


  buf

  (
    g900_n_spl_,
    g900_n
  );


  buf

  (
    g900_p_spl_,
    g900_p
  );


  buf

  (
    g891_n_spl_,
    g891_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    g891_p_spl_,
    g891_p
  );


  buf

  (
    g902_n_spl_,
    g902_n
  );


  buf

  (
    g903_n_spl_,
    g903_n
  );


  buf

  (
    g903_p_spl_,
    g903_p
  );


  buf

  (
    g905_p_spl_,
    g905_p
  );


  buf

  (
    g890_p_spl_,
    g890_p
  );


  buf

  (
    n2821_lo_p_spl_,
    n2821_lo_p
  );


  buf

  (
    n2821_lo_p_spl_0,
    n2821_lo_p_spl_
  );


  buf

  (
    n2821_lo_p_spl_00,
    n2821_lo_p_spl_0
  );


  buf

  (
    n2821_lo_p_spl_000,
    n2821_lo_p_spl_00
  );


  buf

  (
    n2821_lo_p_spl_001,
    n2821_lo_p_spl_00
  );


  buf

  (
    n2821_lo_p_spl_01,
    n2821_lo_p_spl_0
  );


  buf

  (
    n2821_lo_p_spl_1,
    n2821_lo_p_spl_
  );


  buf

  (
    n2821_lo_p_spl_10,
    n2821_lo_p_spl_1
  );


  buf

  (
    n2821_lo_p_spl_11,
    n2821_lo_p_spl_1
  );


  buf

  (
    n2821_lo_n_spl_,
    n2821_lo_n
  );


  buf

  (
    n2821_lo_n_spl_0,
    n2821_lo_n_spl_
  );


  buf

  (
    n2821_lo_n_spl_00,
    n2821_lo_n_spl_0
  );


  buf

  (
    n2821_lo_n_spl_01,
    n2821_lo_n_spl_0
  );


  buf

  (
    n2821_lo_n_spl_1,
    n2821_lo_n_spl_
  );


  buf

  (
    n2821_lo_n_spl_10,
    n2821_lo_n_spl_1
  );


  buf

  (
    n2821_lo_n_spl_11,
    n2821_lo_n_spl_1
  );


  buf

  (
    g839_n_spl_,
    g839_n
  );


  buf

  (
    g789_n_spl_,
    g789_n
  );


  buf

  (
    g739_n_spl_,
    g739_n
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g927_p_spl_,
    g927_p
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g927_n_spl_,
    g927_n
  );


  buf

  (
    g928_p_spl_,
    g928_p
  );


  buf

  (
    g924_n_spl_,
    g924_n
  );


  buf

  (
    g930_p_spl_,
    g930_p
  );


  buf

  (
    g924_p_spl_,
    g924_p
  );


  buf

  (
    g930_n_spl_,
    g930_n
  );


  buf

  (
    g931_p_spl_,
    g931_p
  );


  buf

  (
    g937_n_spl_,
    g937_n
  );


  buf

  (
    g939_p_spl_,
    g939_p
  );


  buf

  (
    g937_p_spl_,
    g937_p
  );


  buf

  (
    g939_n_spl_,
    g939_n
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    g936_n_spl_,
    g936_n
  );


  buf

  (
    g942_p_spl_,
    g942_p
  );


  buf

  (
    g936_p_spl_,
    g936_p
  );


  buf

  (
    g942_n_spl_,
    g942_n
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g949_n_spl_,
    g949_n
  );


  buf

  (
    g951_p_spl_,
    g951_p
  );


  buf

  (
    g949_p_spl_,
    g949_p
  );


  buf

  (
    g951_n_spl_,
    g951_n
  );


  buf

  (
    g952_p_spl_,
    g952_p
  );


  buf

  (
    g948_n_spl_,
    g948_n
  );


  buf

  (
    g954_p_spl_,
    g954_p
  );


  buf

  (
    g948_p_spl_,
    g948_p
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g955_p_spl_,
    g955_p
  );


  buf

  (
    g867_n_spl_,
    g867_n
  );


  buf

  (
    g889_p_spl_,
    g889_p
  );


  buf

  (
    g865_p_spl_,
    g865_p
  );


  buf

  (
    n6025_o2_p_spl_,
    n6025_o2_p
  );


  buf

  (
    n6025_o2_p_spl_0,
    n6025_o2_p_spl_
  );


  buf

  (
    n6025_o2_p_spl_00,
    n6025_o2_p_spl_0
  );


  buf

  (
    n6025_o2_p_spl_01,
    n6025_o2_p_spl_0
  );


  buf

  (
    n6025_o2_p_spl_1,
    n6025_o2_p_spl_
  );


  buf

  (
    n6025_o2_n_spl_,
    n6025_o2_n
  );


  buf

  (
    n6025_o2_n_spl_0,
    n6025_o2_n_spl_
  );


  buf

  (
    n6025_o2_n_spl_00,
    n6025_o2_n_spl_0
  );


  buf

  (
    n6025_o2_n_spl_1,
    n6025_o2_n_spl_
  );


  buf

  (
    n1003_o2_p_spl_,
    n1003_o2_p
  );


  buf

  (
    n1003_o2_n_spl_,
    n1003_o2_n
  );


  buf

  (
    g965_n_spl_,
    g965_n
  );


  buf

  (
    g966_p_spl_,
    g966_p
  );


  buf

  (
    g965_p_spl_,
    g965_p
  );


  buf

  (
    g966_n_spl_,
    g966_n
  );


  buf

  (
    g967_n_spl_,
    g967_n
  );


  buf

  (
    g967_p_spl_,
    g967_p
  );


  buf

  (
    g964_n_spl_,
    g964_n
  );


  buf

  (
    g969_p_spl_,
    g969_p
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g969_n_spl_,
    g969_n
  );


  buf

  (
    g970_n_spl_,
    g970_n
  );


  buf

  (
    g970_p_spl_,
    g970_p
  );


  buf

  (
    g963_n_spl_,
    g963_n
  );


  buf

  (
    g972_p_spl_,
    g972_p
  );


  buf

  (
    g963_p_spl_,
    g963_p
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g973_n_spl_,
    g973_n
  );


  buf

  (
    g973_p_spl_,
    g973_p
  );


  buf

  (
    g962_n_spl_,
    g962_n
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    g962_p_spl_,
    g962_p
  );


  buf

  (
    g975_n_spl_,
    g975_n
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    g976_p_spl_,
    g976_p
  );


  buf

  (
    g961_n_spl_,
    g961_n
  );


  buf

  (
    g978_p_spl_,
    g978_p
  );


  buf

  (
    g961_p_spl_,
    g961_p
  );


  buf

  (
    g978_n_spl_,
    g978_n
  );


  buf

  (
    g979_n_spl_,
    g979_n
  );


  buf

  (
    g979_p_spl_,
    g979_p
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g981_p_spl_,
    g981_p
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g981_n_spl_,
    g981_n
  );


  buf

  (
    g982_n_spl_,
    g982_n
  );


  buf

  (
    g982_p_spl_,
    g982_p
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_01,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_000,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_001,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_01,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_010,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_011,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_10,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_100,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_101,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_11,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_110,
    G17_p_spl_11
  );


  buf

  (
    G17_p_spl_111,
    G17_p_spl_11
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_000,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_001,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_01,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_010,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_011,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_10,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_100,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_101,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_11,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_110,
    G17_n_spl_11
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_000,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_001,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_01,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_010,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_011,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_10,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_100,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_101,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_11,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_110,
    G18_p_spl_11
  );


  buf

  (
    G18_p_spl_111,
    G18_p_spl_11
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_000,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_001,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_01,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_010,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_011,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_10,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_100,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_101,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_11,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_110,
    G18_n_spl_11
  );


  buf

  (
    G18_n_spl_111,
    G18_n_spl_11
  );


  buf

  (
    g984_p_spl_,
    g984_p
  );


  buf

  (
    g907_p_spl_,
    g907_p
  );


  buf

  (
    n2758_lo_p_spl_,
    n2758_lo_p
  );


  buf

  (
    n2758_lo_p_spl_0,
    n2758_lo_p_spl_
  );


  buf

  (
    n2758_lo_p_spl_00,
    n2758_lo_p_spl_0
  );


  buf

  (
    n2758_lo_p_spl_000,
    n2758_lo_p_spl_00
  );


  buf

  (
    n2758_lo_p_spl_001,
    n2758_lo_p_spl_00
  );


  buf

  (
    n2758_lo_p_spl_01,
    n2758_lo_p_spl_0
  );


  buf

  (
    n2758_lo_p_spl_010,
    n2758_lo_p_spl_01
  );


  buf

  (
    n2758_lo_p_spl_011,
    n2758_lo_p_spl_01
  );


  buf

  (
    n2758_lo_p_spl_1,
    n2758_lo_p_spl_
  );


  buf

  (
    n2758_lo_p_spl_10,
    n2758_lo_p_spl_1
  );


  buf

  (
    n2758_lo_p_spl_100,
    n2758_lo_p_spl_10
  );


  buf

  (
    n2758_lo_p_spl_101,
    n2758_lo_p_spl_10
  );


  buf

  (
    n2758_lo_p_spl_11,
    n2758_lo_p_spl_1
  );


  buf

  (
    n2758_lo_n_spl_,
    n2758_lo_n
  );


  buf

  (
    n2758_lo_n_spl_0,
    n2758_lo_n_spl_
  );


  buf

  (
    n2758_lo_n_spl_00,
    n2758_lo_n_spl_0
  );


  buf

  (
    n2758_lo_n_spl_000,
    n2758_lo_n_spl_00
  );


  buf

  (
    n2758_lo_n_spl_001,
    n2758_lo_n_spl_00
  );


  buf

  (
    n2758_lo_n_spl_01,
    n2758_lo_n_spl_0
  );


  buf

  (
    n2758_lo_n_spl_010,
    n2758_lo_n_spl_01
  );


  buf

  (
    n2758_lo_n_spl_011,
    n2758_lo_n_spl_01
  );


  buf

  (
    n2758_lo_n_spl_1,
    n2758_lo_n_spl_
  );


  buf

  (
    n2758_lo_n_spl_10,
    n2758_lo_n_spl_1
  );


  buf

  (
    n2758_lo_n_spl_100,
    n2758_lo_n_spl_10
  );


  buf

  (
    n2758_lo_n_spl_101,
    n2758_lo_n_spl_10
  );


  buf

  (
    n2758_lo_n_spl_11,
    n2758_lo_n_spl_1
  );


  buf

  (
    g985_p_spl_,
    g985_p
  );


  buf

  (
    g986_p_spl_,
    g986_p
  );


  buf

  (
    g906_p_spl_,
    g906_p
  );


  buf

  (
    lo010_buf_o2_p_spl_,
    lo010_buf_o2_p
  );


  buf

  (
    lo010_buf_o2_p_spl_0,
    lo010_buf_o2_p_spl_
  );


  buf

  (
    lo010_buf_o2_p_spl_00,
    lo010_buf_o2_p_spl_0
  );


  buf

  (
    lo010_buf_o2_p_spl_1,
    lo010_buf_o2_p_spl_
  );


  buf

  (
    lo010_buf_o2_n_spl_,
    lo010_buf_o2_n
  );


  buf

  (
    lo010_buf_o2_n_spl_0,
    lo010_buf_o2_n_spl_
  );


  buf

  (
    lo010_buf_o2_n_spl_1,
    lo010_buf_o2_n_spl_
  );


  buf

  (
    n601_o2_n_spl_,
    n601_o2_n
  );


  buf

  (
    n625_o2_p_spl_,
    n625_o2_p
  );


  buf

  (
    n601_o2_p_spl_,
    n601_o2_p
  );


  buf

  (
    n625_o2_n_spl_,
    n625_o2_n
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    g994_n_spl_,
    g994_n
  );


  buf

  (
    g997_p_spl_,
    g997_p
  );


  buf

  (
    g994_p_spl_,
    g994_p
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g998_n_spl_,
    g998_n
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    g993_n_spl_,
    g993_n
  );


  buf

  (
    g1000_p_spl_,
    g1000_p
  );


  buf

  (
    g993_p_spl_,
    g993_p
  );


  buf

  (
    g1000_n_spl_,
    g1000_n
  );


  buf

  (
    g1001_n_spl_,
    g1001_n
  );


  buf

  (
    g1001_p_spl_,
    g1001_p
  );


  buf

  (
    g992_n_spl_,
    g992_n
  );


  buf

  (
    g1003_p_spl_,
    g1003_p
  );


  buf

  (
    g992_p_spl_,
    g992_p
  );


  buf

  (
    g1003_n_spl_,
    g1003_n
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_p_spl_,
    g1004_p
  );


  buf

  (
    g991_n_spl_,
    g991_n
  );


  buf

  (
    g1006_p_spl_,
    g1006_p
  );


  buf

  (
    g991_p_spl_,
    g991_p
  );


  buf

  (
    g1006_n_spl_,
    g1006_n
  );


  buf

  (
    g1007_n_spl_,
    g1007_n
  );


  buf

  (
    g1007_p_spl_,
    g1007_p
  );


  buf

  (
    g990_n_spl_,
    g990_n
  );


  buf

  (
    g1009_p_spl_,
    g1009_p
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g1009_n_spl_,
    g1009_n
  );


  buf

  (
    g1010_n_spl_,
    g1010_n
  );


  buf

  (
    g1010_p_spl_,
    g1010_p
  );


  buf

  (
    g959_p_spl_,
    g959_p
  );


  buf

  (
    g958_n_spl_,
    g958_n
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_000,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_001,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_01,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_010,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_011,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_10,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_100,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_101,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_11,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_110,
    G19_p_spl_11
  );


  buf

  (
    G19_p_spl_111,
    G19_p_spl_11
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_000,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_001,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_01,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_010,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_011,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_10,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_100,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_101,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_11,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_110,
    G19_n_spl_11
  );


  buf

  (
    G19_n_spl_111,
    G19_n_spl_11
  );


  buf

  (
    n1811_o2_n_spl_,
    n1811_o2_n
  );


  buf

  (
    n1811_o2_p_spl_,
    n1811_o2_p
  );


  buf

  (
    n6036_o2_p_spl_,
    n6036_o2_p
  );


  buf

  (
    n6036_o2_p_spl_0,
    n6036_o2_p_spl_
  );


  buf

  (
    n6036_o2_p_spl_00,
    n6036_o2_p_spl_0
  );


  buf

  (
    n6036_o2_p_spl_1,
    n6036_o2_p_spl_
  );


  buf

  (
    lo094_buf_o2_p_spl_,
    lo094_buf_o2_p
  );


  buf

  (
    n6036_o2_n_spl_,
    n6036_o2_n
  );


  buf

  (
    n6036_o2_n_spl_0,
    n6036_o2_n_spl_
  );


  buf

  (
    lo094_buf_o2_n_spl_,
    lo094_buf_o2_n
  );


  buf

  (
    n1889_o2_p_spl_,
    n1889_o2_p
  );


  buf

  (
    n1889_o2_n_spl_,
    n1889_o2_n
  );


  buf

  (
    g1018_n_spl_,
    g1018_n
  );


  buf

  (
    g1019_p_spl_,
    g1019_p
  );


  buf

  (
    g1018_p_spl_,
    g1018_p
  );


  buf

  (
    g1019_n_spl_,
    g1019_n
  );


  buf

  (
    g1020_n_spl_,
    g1020_n
  );


  buf

  (
    g1020_p_spl_,
    g1020_p
  );


  buf

  (
    g1017_n_spl_,
    g1017_n
  );


  buf

  (
    g1022_p_spl_,
    g1022_p
  );


  buf

  (
    g1017_p_spl_,
    g1017_p
  );


  buf

  (
    g1022_n_spl_,
    g1022_n
  );


  buf

  (
    n6035_o2_p_spl_,
    n6035_o2_p
  );


  buf

  (
    n6035_o2_p_spl_0,
    n6035_o2_p_spl_
  );


  buf

  (
    n6035_o2_p_spl_1,
    n6035_o2_p_spl_
  );


  buf

  (
    lo098_buf_o2_p_spl_,
    lo098_buf_o2_p
  );


  buf

  (
    lo098_buf_o2_p_spl_0,
    lo098_buf_o2_p_spl_
  );


  buf

  (
    lo098_buf_o2_p_spl_00,
    lo098_buf_o2_p_spl_0
  );


  buf

  (
    lo098_buf_o2_p_spl_1,
    lo098_buf_o2_p_spl_
  );


  buf

  (
    n6035_o2_n_spl_,
    n6035_o2_n
  );


  buf

  (
    n6035_o2_n_spl_0,
    n6035_o2_n_spl_
  );


  buf

  (
    lo098_buf_o2_n_spl_,
    lo098_buf_o2_n
  );


  buf

  (
    lo098_buf_o2_n_spl_0,
    lo098_buf_o2_n_spl_
  );


  buf

  (
    lo098_buf_o2_n_spl_00,
    lo098_buf_o2_n_spl_0
  );


  buf

  (
    lo098_buf_o2_n_spl_1,
    lo098_buf_o2_n_spl_
  );


  buf

  (
    g1023_n_spl_,
    g1023_n
  );


  buf

  (
    g1023_p_spl_,
    g1023_p
  );


  buf

  (
    g1024_n_spl_,
    g1024_n
  );


  buf

  (
    g1026_p_spl_,
    g1026_p
  );


  buf

  (
    g1024_p_spl_,
    g1024_p
  );


  buf

  (
    g1026_n_spl_,
    g1026_n
  );


  buf

  (
    g1027_n_spl_,
    g1027_n
  );


  buf

  (
    g1027_p_spl_,
    g1027_p
  );


  buf

  (
    n6037_o2_p_spl_,
    n6037_o2_p
  );


  buf

  (
    n6037_o2_p_spl_0,
    n6037_o2_p_spl_
  );


  buf

  (
    n6037_o2_p_spl_1,
    n6037_o2_p_spl_
  );


  buf

  (
    n6037_o2_n_spl_,
    n6037_o2_n
  );


  buf

  (
    n6037_o2_n_spl_0,
    n6037_o2_n_spl_
  );


  buf

  (
    g1030_n_spl_,
    g1030_n
  );


  buf

  (
    g1031_n_spl_,
    g1031_n
  );


  buf

  (
    g1030_p_spl_,
    g1030_p
  );


  buf

  (
    g1031_p_spl_,
    g1031_p
  );


  buf

  (
    g1032_n_spl_,
    g1032_n
  );


  buf

  (
    g1032_p_spl_,
    g1032_p
  );


  buf

  (
    g1029_n_spl_,
    g1029_n
  );


  buf

  (
    g1034_p_spl_,
    g1034_p
  );


  buf

  (
    g1029_p_spl_,
    g1029_p
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    g1035_n_spl_,
    g1035_n
  );


  buf

  (
    g1035_p_spl_,
    g1035_p
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    g1037_p_spl_,
    g1037_p
  );


  buf

  (
    g1028_p_spl_,
    g1028_p
  );


  buf

  (
    g1037_n_spl_,
    g1037_n
  );


  buf

  (
    g1038_n_spl_,
    g1038_n
  );


  buf

  (
    g1038_p_spl_,
    g1038_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1041_p_spl_,
    g1041_p
  );


  buf

  (
    g1039_p_spl_,
    g1039_p
  );


  buf

  (
    g1041_n_spl_,
    g1041_n
  );


  buf

  (
    g1042_n_spl_,
    g1042_n
  );


  buf

  (
    g1042_p_spl_,
    g1042_p
  );


  buf

  (
    g1045_n_spl_,
    g1045_n
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1045_p_spl_,
    g1045_p
  );


  buf

  (
    g1046_p_spl_,
    g1046_p
  );


  buf

  (
    g1047_n_spl_,
    g1047_n
  );


  buf

  (
    g1047_p_spl_,
    g1047_p
  );


  buf

  (
    g1044_n_spl_,
    g1044_n
  );


  buf

  (
    g1049_p_spl_,
    g1049_p
  );


  buf

  (
    g1044_p_spl_,
    g1044_p
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1050_n_spl_,
    g1050_n
  );


  buf

  (
    g1050_p_spl_,
    g1050_p
  );


  buf

  (
    g1043_n_spl_,
    g1043_n
  );


  buf

  (
    g1052_p_spl_,
    g1052_p
  );


  buf

  (
    g1043_p_spl_,
    g1043_p
  );


  buf

  (
    g1052_n_spl_,
    g1052_n
  );


  buf

  (
    n1631_o2_n_spl_,
    n1631_o2_n
  );


  buf

  (
    n1631_o2_p_spl_,
    n1631_o2_p
  );


  buf

  (
    n6033_o2_p_spl_,
    n6033_o2_p
  );


  buf

  (
    n6033_o2_p_spl_0,
    n6033_o2_p_spl_
  );


  buf

  (
    n6033_o2_p_spl_00,
    n6033_o2_p_spl_0
  );


  buf

  (
    n6033_o2_p_spl_1,
    n6033_o2_p_spl_
  );


  buf

  (
    n6033_o2_n_spl_,
    n6033_o2_n
  );


  buf

  (
    n6033_o2_n_spl_0,
    n6033_o2_n_spl_
  );


  buf

  (
    n1725_o2_p_spl_,
    n1725_o2_p
  );


  buf

  (
    n1725_o2_n_spl_,
    n1725_o2_n
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1056_p_spl_,
    g1056_p
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    g1056_n_spl_,
    g1056_n
  );


  buf

  (
    g1057_n_spl_,
    g1057_n
  );


  buf

  (
    g1057_p_spl_,
    g1057_p
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g1059_p_spl_,
    g1059_p
  );


  buf

  (
    g1054_p_spl_,
    g1054_p
  );


  buf

  (
    g1059_n_spl_,
    g1059_n
  );


  buf

  (
    n6032_o2_p_spl_,
    n6032_o2_p
  );


  buf

  (
    n6032_o2_p_spl_0,
    n6032_o2_p_spl_
  );


  buf

  (
    n6032_o2_p_spl_1,
    n6032_o2_p_spl_
  );


  buf

  (
    n6032_o2_n_spl_,
    n6032_o2_n
  );


  buf

  (
    n6032_o2_n_spl_0,
    n6032_o2_n_spl_
  );


  buf

  (
    g1060_n_spl_,
    g1060_n
  );


  buf

  (
    g1060_p_spl_,
    g1060_p
  );


  buf

  (
    g1061_n_spl_,
    g1061_n
  );


  buf

  (
    g1063_p_spl_,
    g1063_p
  );


  buf

  (
    g1061_p_spl_,
    g1061_p
  );


  buf

  (
    g1063_n_spl_,
    g1063_n
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1064_p_spl_,
    g1064_p
  );


  buf

  (
    n6034_o2_p_spl_,
    n6034_o2_p
  );


  buf

  (
    n6034_o2_p_spl_0,
    n6034_o2_p_spl_
  );


  buf

  (
    n6034_o2_p_spl_1,
    n6034_o2_p_spl_
  );


  buf

  (
    n6034_o2_n_spl_,
    n6034_o2_n
  );


  buf

  (
    n6034_o2_n_spl_0,
    n6034_o2_n_spl_
  );


  buf

  (
    g1069_n_spl_,
    g1069_n
  );


  buf

  (
    g1070_p_spl_,
    g1070_p
  );


  buf

  (
    g1069_p_spl_,
    g1069_p
  );


  buf

  (
    g1070_n_spl_,
    g1070_n
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1071_p_spl_,
    g1071_p
  );


  buf

  (
    g1068_n_spl_,
    g1068_n
  );


  buf

  (
    g1073_p_spl_,
    g1073_p
  );


  buf

  (
    g1068_p_spl_,
    g1068_p
  );


  buf

  (
    g1073_n_spl_,
    g1073_n
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g1074_p_spl_,
    g1074_p
  );


  buf

  (
    g1067_n_spl_,
    g1067_n
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1067_p_spl_,
    g1067_p
  );


  buf

  (
    g1076_n_spl_,
    g1076_n
  );


  buf

  (
    g1077_n_spl_,
    g1077_n
  );


  buf

  (
    g1077_p_spl_,
    g1077_p
  );


  buf

  (
    g1066_n_spl_,
    g1066_n
  );


  buf

  (
    g1079_p_spl_,
    g1079_p
  );


  buf

  (
    g1066_p_spl_,
    g1066_p
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1080_n_spl_,
    g1080_n
  );


  buf

  (
    g1080_p_spl_,
    g1080_p
  );


  buf

  (
    g1065_n_spl_,
    g1065_n
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1065_p_spl_,
    g1065_p
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    g1083_n_spl_,
    g1083_n
  );


  buf

  (
    g1083_p_spl_,
    g1083_p
  );


  buf

  (
    g1084_n_spl_,
    g1084_n
  );


  buf

  (
    g1086_p_spl_,
    g1086_p
  );


  buf

  (
    g1084_p_spl_,
    g1084_p
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g1087_n_spl_,
    g1087_n
  );


  buf

  (
    g1087_p_spl_,
    g1087_p
  );


  buf

  (
    g1092_n_spl_,
    g1092_n
  );


  buf

  (
    g1094_p_spl_,
    g1094_p
  );


  buf

  (
    g1092_p_spl_,
    g1092_p
  );


  buf

  (
    g1094_n_spl_,
    g1094_n
  );


  buf

  (
    g1095_n_spl_,
    g1095_n
  );


  buf

  (
    g1095_p_spl_,
    g1095_p
  );


  buf

  (
    g1091_n_spl_,
    g1091_n
  );


  buf

  (
    g1097_p_spl_,
    g1097_p
  );


  buf

  (
    g1091_p_spl_,
    g1091_p
  );


  buf

  (
    g1097_n_spl_,
    g1097_n
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    g1098_p_spl_,
    g1098_p
  );


  buf

  (
    g1090_n_spl_,
    g1090_n
  );


  buf

  (
    g1100_p_spl_,
    g1100_p
  );


  buf

  (
    g1090_p_spl_,
    g1090_p
  );


  buf

  (
    g1100_n_spl_,
    g1100_n
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    g1101_p_spl_,
    g1101_p
  );


  buf

  (
    g1089_n_spl_,
    g1089_n
  );


  buf

  (
    g1103_p_spl_,
    g1103_p
  );


  buf

  (
    g1089_p_spl_,
    g1089_p
  );


  buf

  (
    g1103_n_spl_,
    g1103_n
  );


  buf

  (
    g1104_n_spl_,
    g1104_n
  );


  buf

  (
    g1104_p_spl_,
    g1104_p
  );


  buf

  (
    g1088_n_spl_,
    g1088_n
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g1106_n_spl_,
    g1106_n
  );


  buf

  (
    n6029_o2_p_spl_,
    n6029_o2_p
  );


  buf

  (
    n6029_o2_p_spl_0,
    n6029_o2_p_spl_
  );


  buf

  (
    n6029_o2_p_spl_00,
    n6029_o2_p_spl_0
  );


  buf

  (
    n6029_o2_p_spl_1,
    n6029_o2_p_spl_
  );


  buf

  (
    n6029_o2_n_spl_,
    n6029_o2_n
  );


  buf

  (
    n6029_o2_n_spl_0,
    n6029_o2_n_spl_
  );


  buf

  (
    n6029_o2_n_spl_1,
    n6029_o2_n_spl_
  );


  buf

  (
    n1420_o2_p_spl_,
    n1420_o2_p
  );


  buf

  (
    n1420_o2_n_spl_,
    n1420_o2_n
  );


  buf

  (
    g1108_n_spl_,
    g1108_n
  );


  buf

  (
    g1109_p_spl_,
    g1109_p
  );


  buf

  (
    g1108_p_spl_,
    g1108_p
  );


  buf

  (
    g1109_n_spl_,
    g1109_n
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1110_p_spl_,
    g1110_p
  );


  buf

  (
    n6030_o2_p_spl_,
    n6030_o2_p
  );


  buf

  (
    n6030_o2_p_spl_0,
    n6030_o2_p_spl_
  );


  buf

  (
    n6030_o2_p_spl_00,
    n6030_o2_p_spl_0
  );


  buf

  (
    n6030_o2_p_spl_1,
    n6030_o2_p_spl_
  );


  buf

  (
    n6030_o2_n_spl_,
    n6030_o2_n
  );


  buf

  (
    n6030_o2_n_spl_0,
    n6030_o2_n_spl_
  );


  buf

  (
    n1529_o2_p_spl_,
    n1529_o2_p
  );


  buf

  (
    n1529_o2_n_spl_,
    n1529_o2_n
  );


  buf

  (
    g1112_n_spl_,
    g1112_n
  );


  buf

  (
    g1113_p_spl_,
    g1113_p
  );


  buf

  (
    g1112_p_spl_,
    g1112_p
  );


  buf

  (
    g1113_n_spl_,
    g1113_n
  );


  buf

  (
    g1114_n_spl_,
    g1114_n
  );


  buf

  (
    g1114_p_spl_,
    g1114_p
  );


  buf

  (
    g1111_n_spl_,
    g1111_n
  );


  buf

  (
    g1116_p_spl_,
    g1116_p
  );


  buf

  (
    g1111_p_spl_,
    g1111_p
  );


  buf

  (
    g1116_n_spl_,
    g1116_n
  );


  buf

  (
    g1117_n_spl_,
    g1117_n
  );


  buf

  (
    g1117_p_spl_,
    g1117_p
  );


  buf

  (
    g1118_n_spl_,
    g1118_n
  );


  buf

  (
    g1120_p_spl_,
    g1120_p
  );


  buf

  (
    g1118_p_spl_,
    g1118_p
  );


  buf

  (
    g1120_n_spl_,
    g1120_n
  );


  buf

  (
    g1121_n_spl_,
    g1121_n
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    n6031_o2_p_spl_,
    n6031_o2_p
  );


  buf

  (
    n6031_o2_p_spl_0,
    n6031_o2_p_spl_
  );


  buf

  (
    n6031_o2_p_spl_1,
    n6031_o2_p_spl_
  );


  buf

  (
    n6031_o2_n_spl_,
    n6031_o2_n
  );


  buf

  (
    n6031_o2_n_spl_0,
    n6031_o2_n_spl_
  );


  buf

  (
    g1126_n_spl_,
    g1126_n
  );


  buf

  (
    g1127_p_spl_,
    g1127_p
  );


  buf

  (
    g1126_p_spl_,
    g1126_p
  );


  buf

  (
    g1127_n_spl_,
    g1127_n
  );


  buf

  (
    g1128_n_spl_,
    g1128_n
  );


  buf

  (
    g1128_p_spl_,
    g1128_p
  );


  buf

  (
    g1125_n_spl_,
    g1125_n
  );


  buf

  (
    g1130_p_spl_,
    g1130_p
  );


  buf

  (
    g1125_p_spl_,
    g1125_p
  );


  buf

  (
    g1130_n_spl_,
    g1130_n
  );


  buf

  (
    g1131_n_spl_,
    g1131_n
  );


  buf

  (
    g1131_p_spl_,
    g1131_p
  );


  buf

  (
    g1124_n_spl_,
    g1124_n
  );


  buf

  (
    g1133_p_spl_,
    g1133_p
  );


  buf

  (
    g1124_p_spl_,
    g1124_p
  );


  buf

  (
    g1133_n_spl_,
    g1133_n
  );


  buf

  (
    g1134_n_spl_,
    g1134_n
  );


  buf

  (
    g1134_p_spl_,
    g1134_p
  );


  buf

  (
    g1123_n_spl_,
    g1123_n
  );


  buf

  (
    g1136_p_spl_,
    g1136_p
  );


  buf

  (
    g1123_p_spl_,
    g1123_p
  );


  buf

  (
    g1136_n_spl_,
    g1136_n
  );


  buf

  (
    g1137_n_spl_,
    g1137_n
  );


  buf

  (
    g1137_p_spl_,
    g1137_p
  );


  buf

  (
    g1122_n_spl_,
    g1122_n
  );


  buf

  (
    g1139_p_spl_,
    g1139_p
  );


  buf

  (
    g1122_p_spl_,
    g1122_p
  );


  buf

  (
    g1139_n_spl_,
    g1139_n
  );


  buf

  (
    g1140_n_spl_,
    g1140_n
  );


  buf

  (
    g1140_p_spl_,
    g1140_p
  );


  buf

  (
    g1141_n_spl_,
    g1141_n
  );


  buf

  (
    g1143_p_spl_,
    g1143_p
  );


  buf

  (
    g1141_p_spl_,
    g1141_p
  );


  buf

  (
    g1143_n_spl_,
    g1143_n
  );


  buf

  (
    g1144_n_spl_,
    g1144_n
  );


  buf

  (
    g1144_p_spl_,
    g1144_p
  );


  buf

  (
    g1149_n_spl_,
    g1149_n
  );


  buf

  (
    g1151_p_spl_,
    g1151_p
  );


  buf

  (
    g1149_p_spl_,
    g1149_p
  );


  buf

  (
    g1151_n_spl_,
    g1151_n
  );


  buf

  (
    g1152_n_spl_,
    g1152_n
  );


  buf

  (
    g1152_p_spl_,
    g1152_p
  );


  buf

  (
    g1148_n_spl_,
    g1148_n
  );


  buf

  (
    g1154_p_spl_,
    g1154_p
  );


  buf

  (
    g1148_p_spl_,
    g1148_p
  );


  buf

  (
    g1154_n_spl_,
    g1154_n
  );


  buf

  (
    g1155_n_spl_,
    g1155_n
  );


  buf

  (
    g1155_p_spl_,
    g1155_p
  );


  buf

  (
    g1147_n_spl_,
    g1147_n
  );


  buf

  (
    g1157_p_spl_,
    g1157_p
  );


  buf

  (
    g1147_p_spl_,
    g1147_p
  );


  buf

  (
    g1157_n_spl_,
    g1157_n
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1158_p_spl_,
    g1158_p
  );


  buf

  (
    g1146_n_spl_,
    g1146_n
  );


  buf

  (
    g1160_p_spl_,
    g1160_p
  );


  buf

  (
    g1146_p_spl_,
    g1146_p
  );


  buf

  (
    g1160_n_spl_,
    g1160_n
  );


  buf

  (
    g1161_n_spl_,
    g1161_n
  );


  buf

  (
    g1161_p_spl_,
    g1161_p
  );


  buf

  (
    g1145_n_spl_,
    g1145_n
  );


  buf

  (
    g1163_p_spl_,
    g1163_p
  );


  buf

  (
    g1145_p_spl_,
    g1145_p
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    n6026_o2_p_spl_,
    n6026_o2_p
  );


  buf

  (
    n6026_o2_p_spl_0,
    n6026_o2_p_spl_
  );


  buf

  (
    n6026_o2_p_spl_00,
    n6026_o2_p_spl_0
  );


  buf

  (
    n6026_o2_p_spl_01,
    n6026_o2_p_spl_0
  );


  buf

  (
    n6026_o2_p_spl_1,
    n6026_o2_p_spl_
  );


  buf

  (
    n6026_o2_n_spl_,
    n6026_o2_n
  );


  buf

  (
    n6026_o2_n_spl_0,
    n6026_o2_n_spl_
  );


  buf

  (
    n6026_o2_n_spl_00,
    n6026_o2_n_spl_0
  );


  buf

  (
    n6026_o2_n_spl_1,
    n6026_o2_n_spl_
  );


  buf

  (
    n1097_o2_p_spl_,
    n1097_o2_p
  );


  buf

  (
    n1097_o2_n_spl_,
    n1097_o2_n
  );


  buf

  (
    g1165_n_spl_,
    g1165_n
  );


  buf

  (
    g1166_p_spl_,
    g1166_p
  );


  buf

  (
    g1165_p_spl_,
    g1165_p
  );


  buf

  (
    g1166_n_spl_,
    g1166_n
  );


  buf

  (
    g1167_n_spl_,
    g1167_n
  );


  buf

  (
    g1167_p_spl_,
    g1167_p
  );


  buf

  (
    n6027_o2_p_spl_,
    n6027_o2_p
  );


  buf

  (
    n6027_o2_p_spl_0,
    n6027_o2_p_spl_
  );


  buf

  (
    n6027_o2_p_spl_00,
    n6027_o2_p_spl_0
  );


  buf

  (
    n6027_o2_p_spl_01,
    n6027_o2_p_spl_0
  );


  buf

  (
    n6027_o2_p_spl_1,
    n6027_o2_p_spl_
  );


  buf

  (
    n6027_o2_n_spl_,
    n6027_o2_n
  );


  buf

  (
    n6027_o2_n_spl_0,
    n6027_o2_n_spl_
  );


  buf

  (
    n6027_o2_n_spl_1,
    n6027_o2_n_spl_
  );


  buf

  (
    n1199_o2_p_spl_,
    n1199_o2_p
  );


  buf

  (
    n1199_o2_n_spl_,
    n1199_o2_n
  );


  buf

  (
    g1169_n_spl_,
    g1169_n
  );


  buf

  (
    g1170_p_spl_,
    g1170_p
  );


  buf

  (
    g1169_p_spl_,
    g1169_p
  );


  buf

  (
    g1170_n_spl_,
    g1170_n
  );


  buf

  (
    g1171_n_spl_,
    g1171_n
  );


  buf

  (
    g1171_p_spl_,
    g1171_p
  );


  buf

  (
    g1168_n_spl_,
    g1168_n
  );


  buf

  (
    g1173_p_spl_,
    g1173_p
  );


  buf

  (
    g1168_p_spl_,
    g1168_p
  );


  buf

  (
    g1173_n_spl_,
    g1173_n
  );


  buf

  (
    g1174_n_spl_,
    g1174_n
  );


  buf

  (
    g1174_p_spl_,
    g1174_p
  );


  buf

  (
    g1175_n_spl_,
    g1175_n
  );


  buf

  (
    g1177_p_spl_,
    g1177_p
  );


  buf

  (
    g1175_p_spl_,
    g1175_p
  );


  buf

  (
    g1177_n_spl_,
    g1177_n
  );


  buf

  (
    g1178_n_spl_,
    g1178_n
  );


  buf

  (
    g1178_p_spl_,
    g1178_p
  );


  buf

  (
    n6028_o2_p_spl_,
    n6028_o2_p
  );


  buf

  (
    n6028_o2_p_spl_0,
    n6028_o2_p_spl_
  );


  buf

  (
    n6028_o2_p_spl_00,
    n6028_o2_p_spl_0
  );


  buf

  (
    n6028_o2_p_spl_1,
    n6028_o2_p_spl_
  );


  buf

  (
    n6028_o2_n_spl_,
    n6028_o2_n
  );


  buf

  (
    n6028_o2_n_spl_0,
    n6028_o2_n_spl_
  );


  buf

  (
    n6028_o2_n_spl_1,
    n6028_o2_n_spl_
  );


  buf

  (
    n1309_o2_p_spl_,
    n1309_o2_p
  );


  buf

  (
    n1309_o2_n_spl_,
    n1309_o2_n
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1183_p_spl_,
    g1183_p
  );


  buf

  (
    g1182_p_spl_,
    g1182_p
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1184_n_spl_,
    g1184_n
  );


  buf

  (
    g1184_p_spl_,
    g1184_p
  );


  buf

  (
    g1181_n_spl_,
    g1181_n
  );


  buf

  (
    g1186_p_spl_,
    g1186_p
  );


  buf

  (
    g1181_p_spl_,
    g1181_p
  );


  buf

  (
    g1186_n_spl_,
    g1186_n
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1187_p_spl_,
    g1187_p
  );


  buf

  (
    g1180_n_spl_,
    g1180_n
  );


  buf

  (
    g1189_p_spl_,
    g1189_p
  );


  buf

  (
    g1180_p_spl_,
    g1180_p
  );


  buf

  (
    g1189_n_spl_,
    g1189_n
  );


  buf

  (
    g1190_n_spl_,
    g1190_n
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1179_n_spl_,
    g1179_n
  );


  buf

  (
    g1192_p_spl_,
    g1192_p
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g1192_n_spl_,
    g1192_n
  );


  buf

  (
    g1193_n_spl_,
    g1193_n
  );


  buf

  (
    g1193_p_spl_,
    g1193_p
  );


  buf

  (
    g1194_n_spl_,
    g1194_n
  );


  buf

  (
    g1196_p_spl_,
    g1196_p
  );


  buf

  (
    g1194_p_spl_,
    g1194_p
  );


  buf

  (
    g1196_n_spl_,
    g1196_n
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1197_p_spl_,
    g1197_p
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1204_p_spl_,
    g1204_p
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1204_n_spl_,
    g1204_n
  );


  buf

  (
    g1205_n_spl_,
    g1205_n
  );


  buf

  (
    g1205_p_spl_,
    g1205_p
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    g1207_p_spl_,
    g1207_p
  );


  buf

  (
    g1201_p_spl_,
    g1201_p
  );


  buf

  (
    g1207_n_spl_,
    g1207_n
  );


  buf

  (
    g1208_n_spl_,
    g1208_n
  );


  buf

  (
    g1208_p_spl_,
    g1208_p
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1210_p_spl_,
    g1210_p
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1210_n_spl_,
    g1210_n
  );


  buf

  (
    g1211_n_spl_,
    g1211_n
  );


  buf

  (
    g1211_p_spl_,
    g1211_p
  );


  buf

  (
    g1199_n_spl_,
    g1199_n
  );


  buf

  (
    g1213_p_spl_,
    g1213_p
  );


  buf

  (
    g1199_p_spl_,
    g1199_p
  );


  buf

  (
    g1213_n_spl_,
    g1213_n
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1198_n_spl_,
    g1198_n
  );


  buf

  (
    g1216_p_spl_,
    g1216_p
  );


  buf

  (
    g1198_p_spl_,
    g1198_p
  );


  buf

  (
    g1216_n_spl_,
    g1216_n
  );


  buf

  (
    g1217_n_spl_,
    g1217_n
  );


  buf

  (
    g1217_p_spl_,
    g1217_p
  );


  buf

  (
    g1218_n_spl_,
    g1218_n
  );


  buf

  (
    g1220_p_spl_,
    g1220_p
  );


  buf

  (
    g1218_p_spl_,
    g1218_p
  );


  buf

  (
    g1220_n_spl_,
    g1220_n
  );


  buf

  (
    g1221_n_spl_,
    g1221_n
  );


  buf

  (
    g1221_p_spl_,
    g1221_p
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1228_p_spl_,
    g1228_p
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1228_n_spl_,
    g1228_n
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1225_n_spl_,
    g1225_n
  );


  buf

  (
    g1231_p_spl_,
    g1231_p
  );


  buf

  (
    g1225_p_spl_,
    g1225_p
  );


  buf

  (
    g1231_n_spl_,
    g1231_n
  );


  buf

  (
    g1232_n_spl_,
    g1232_n
  );


  buf

  (
    g1232_p_spl_,
    g1232_p
  );


  buf

  (
    g1224_n_spl_,
    g1224_n
  );


  buf

  (
    g1234_p_spl_,
    g1234_p
  );


  buf

  (
    g1224_p_spl_,
    g1224_p
  );


  buf

  (
    g1234_n_spl_,
    g1234_n
  );


  buf

  (
    g1235_n_spl_,
    g1235_n
  );


  buf

  (
    g1235_p_spl_,
    g1235_p
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1237_p_spl_,
    g1237_p
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1237_n_spl_,
    g1237_n
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1222_n_spl_,
    g1222_n
  );


  buf

  (
    g1240_p_spl_,
    g1240_p
  );


  buf

  (
    g1222_p_spl_,
    g1222_p
  );


  buf

  (
    g1240_n_spl_,
    g1240_n
  );


  buf

  (
    g1012_p_spl_,
    g1012_p
  );


  buf

  (
    g988_p_spl_,
    g988_p
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_01,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    g1243_p_spl_,
    g1243_p
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1243_n_spl_,
    g1243_n
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1245_n_spl_,
    g1245_n
  );


  buf

  (
    g1245_n_spl_0,
    g1245_n_spl_
  );


  buf

  (
    g1245_p_spl_,
    g1245_p
  );


  buf

  (
    g1245_p_spl_0,
    g1245_p_spl_
  );


  buf

  (
    g989_n_spl_,
    g989_n
  );


  buf

  (
    g1247_n_spl_,
    g1247_n
  );


  buf

  (
    g989_p_spl_,
    g989_p
  );


  buf

  (
    g989_p_spl_0,
    g989_p_spl_
  );


  buf

  (
    g1247_p_spl_,
    g1247_p
  );


  buf

  (
    g1248_n_spl_,
    g1248_n
  );


  buf

  (
    g1248_p_spl_,
    g1248_p
  );


  buf

  (
    g987_p_spl_,
    g987_p
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    g1259_p_spl_,
    g1259_p
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1259_n_spl_,
    g1259_n
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1256_n_spl_,
    g1256_n
  );


  buf

  (
    g1262_p_spl_,
    g1262_p
  );


  buf

  (
    g1256_p_spl_,
    g1256_p
  );


  buf

  (
    g1262_n_spl_,
    g1262_n
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1255_n_spl_,
    g1255_n
  );


  buf

  (
    g1265_p_spl_,
    g1265_p
  );


  buf

  (
    g1255_p_spl_,
    g1255_p
  );


  buf

  (
    g1265_n_spl_,
    g1265_n
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1269_n_spl_,
    g1269_n
  );


  buf

  (
    g1269_p_spl_,
    g1269_p
  );


  buf

  (
    g1253_n_spl_,
    g1253_n
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1253_p_spl_,
    g1253_p
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1272_n_spl_,
    g1272_n
  );


  buf

  (
    g1272_p_spl_,
    g1272_p
  );


  buf

  (
    g1252_n_spl_,
    g1252_n
  );


  buf

  (
    g1274_p_spl_,
    g1274_p
  );


  buf

  (
    g1252_p_spl_,
    g1252_p
  );


  buf

  (
    g1274_n_spl_,
    g1274_n
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    n1374_o2_n_spl_,
    n1374_o2_n
  );


  buf

  (
    n1392_o2_p_spl_,
    n1392_o2_p
  );


  buf

  (
    n1374_o2_p_spl_,
    n1374_o2_p
  );


  buf

  (
    n1392_o2_n_spl_,
    n1392_o2_n
  );


  buf

  (
    g1279_n_spl_,
    g1279_n
  );


  buf

  (
    g1279_p_spl_,
    g1279_p
  );


  buf

  (
    n1488_o2_n_spl_,
    n1488_o2_n
  );


  buf

  (
    n1501_o2_p_spl_,
    n1501_o2_p
  );


  buf

  (
    n1488_o2_p_spl_,
    n1488_o2_p
  );


  buf

  (
    n1501_o2_n_spl_,
    n1501_o2_n
  );


  buf

  (
    g1281_n_spl_,
    g1281_n
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1280_n_spl_,
    g1280_n
  );


  buf

  (
    g1283_p_spl_,
    g1283_p
  );


  buf

  (
    g1280_p_spl_,
    g1280_p
  );


  buf

  (
    g1283_n_spl_,
    g1283_n
  );


  buf

  (
    lo050_buf_o2_p_spl_,
    lo050_buf_o2_p
  );


  buf

  (
    lo050_buf_o2_p_spl_0,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    lo050_buf_o2_p_spl_1,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    lo050_buf_o2_n_spl_,
    lo050_buf_o2_n
  );


  buf

  (
    lo050_buf_o2_n_spl_0,
    lo050_buf_o2_n_spl_
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1285_n_spl_,
    g1285_n
  );


  buf

  (
    g1287_p_spl_,
    g1287_p
  );


  buf

  (
    g1285_p_spl_,
    g1285_p
  );


  buf

  (
    g1287_n_spl_,
    g1287_n
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    lo054_buf_o2_p_spl_,
    lo054_buf_o2_p
  );


  buf

  (
    lo054_buf_o2_p_spl_0,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    lo054_buf_o2_n_spl_,
    lo054_buf_o2_n
  );


  buf

  (
    lo054_buf_o2_n_spl_0,
    lo054_buf_o2_n_spl_
  );


  buf

  (
    lo058_buf_o2_p_spl_,
    lo058_buf_o2_p
  );


  buf

  (
    lo058_buf_o2_p_spl_0,
    lo058_buf_o2_p_spl_
  );


  buf

  (
    lo058_buf_o2_p_spl_1,
    lo058_buf_o2_p_spl_
  );


  buf

  (
    lo058_buf_o2_n_spl_,
    lo058_buf_o2_n
  );


  buf

  (
    lo058_buf_o2_n_spl_0,
    lo058_buf_o2_n_spl_
  );


  buf

  (
    n1602_o2_n_spl_,
    n1602_o2_n
  );


  buf

  (
    n1603_o2_n_spl_,
    n1603_o2_n
  );


  buf

  (
    n1602_o2_p_spl_,
    n1602_o2_p
  );


  buf

  (
    n1603_o2_p_spl_,
    n1603_o2_p
  );


  buf

  (
    g1293_n_spl_,
    g1293_n
  );


  buf

  (
    g1293_p_spl_,
    g1293_p
  );


  buf

  (
    g1292_n_spl_,
    g1292_n
  );


  buf

  (
    g1295_p_spl_,
    g1295_p
  );


  buf

  (
    g1292_p_spl_,
    g1292_p
  );


  buf

  (
    g1295_n_spl_,
    g1295_n
  );


  buf

  (
    g1296_n_spl_,
    g1296_n
  );


  buf

  (
    g1296_p_spl_,
    g1296_p
  );


  buf

  (
    g1291_n_spl_,
    g1291_n
  );


  buf

  (
    g1298_p_spl_,
    g1298_p
  );


  buf

  (
    g1291_p_spl_,
    g1291_p
  );


  buf

  (
    g1298_n_spl_,
    g1298_n
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1290_n_spl_,
    g1290_n
  );


  buf

  (
    g1301_p_spl_,
    g1301_p
  );


  buf

  (
    g1290_p_spl_,
    g1290_p
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1302_n_spl_,
    g1302_n
  );


  buf

  (
    g1302_p_spl_,
    g1302_p
  );


  buf

  (
    g1289_n_spl_,
    g1289_n
  );


  buf

  (
    g1304_p_spl_,
    g1304_p
  );


  buf

  (
    g1289_p_spl_,
    g1289_p
  );


  buf

  (
    g1304_n_spl_,
    g1304_n
  );


  buf

  (
    g1305_n_spl_,
    g1305_n
  );


  buf

  (
    g1305_p_spl_,
    g1305_p
  );


  buf

  (
    g1306_n_spl_,
    g1306_n
  );


  buf

  (
    g1308_p_spl_,
    g1308_p
  );


  buf

  (
    g1306_p_spl_,
    g1306_p
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1309_n_spl_,
    g1309_n
  );


  buf

  (
    g1309_p_spl_,
    g1309_p
  );


  buf

  (
    lo062_buf_o2_p_spl_,
    lo062_buf_o2_p
  );


  buf

  (
    lo062_buf_o2_p_spl_0,
    lo062_buf_o2_p_spl_
  );


  buf

  (
    lo062_buf_o2_n_spl_,
    lo062_buf_o2_n
  );


  buf

  (
    lo062_buf_o2_n_spl_0,
    lo062_buf_o2_n_spl_
  );


  buf

  (
    g1314_n_spl_,
    g1314_n
  );


  buf

  (
    g1315_n_spl_,
    g1315_n
  );


  buf

  (
    g1314_p_spl_,
    g1314_p
  );


  buf

  (
    g1315_p_spl_,
    g1315_p
  );


  buf

  (
    g1316_n_spl_,
    g1316_n
  );


  buf

  (
    g1316_p_spl_,
    g1316_p
  );


  buf

  (
    g1313_n_spl_,
    g1313_n
  );


  buf

  (
    g1318_p_spl_,
    g1318_p
  );


  buf

  (
    g1313_p_spl_,
    g1313_p
  );


  buf

  (
    g1318_n_spl_,
    g1318_n
  );


  buf

  (
    g1319_n_spl_,
    g1319_n
  );


  buf

  (
    g1319_p_spl_,
    g1319_p
  );


  buf

  (
    g1312_n_spl_,
    g1312_n
  );


  buf

  (
    g1321_p_spl_,
    g1321_p
  );


  buf

  (
    g1312_p_spl_,
    g1312_p
  );


  buf

  (
    g1321_n_spl_,
    g1321_n
  );


  buf

  (
    g1322_n_spl_,
    g1322_n
  );


  buf

  (
    g1322_p_spl_,
    g1322_p
  );


  buf

  (
    g1311_n_spl_,
    g1311_n
  );


  buf

  (
    g1324_p_spl_,
    g1324_p
  );


  buf

  (
    g1311_p_spl_,
    g1311_p
  );


  buf

  (
    g1324_n_spl_,
    g1324_n
  );


  buf

  (
    g1325_n_spl_,
    g1325_n
  );


  buf

  (
    g1325_p_spl_,
    g1325_p
  );


  buf

  (
    g1310_n_spl_,
    g1310_n
  );


  buf

  (
    g1327_p_spl_,
    g1327_p
  );


  buf

  (
    g1310_p_spl_,
    g1310_p
  );


  buf

  (
    g1327_n_spl_,
    g1327_n
  );


  buf

  (
    n1045_o2_n_spl_,
    n1045_o2_n
  );


  buf

  (
    n1069_o2_p_spl_,
    n1069_o2_p
  );


  buf

  (
    n1045_o2_p_spl_,
    n1045_o2_p
  );


  buf

  (
    n1069_o2_n_spl_,
    n1069_o2_n
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    n1147_o2_n_spl_,
    n1147_o2_n
  );


  buf

  (
    n1171_o2_p_spl_,
    n1171_o2_p
  );


  buf

  (
    n1147_o2_p_spl_,
    n1147_o2_p
  );


  buf

  (
    n1171_o2_n_spl_,
    n1171_o2_n
  );


  buf

  (
    g1331_n_spl_,
    g1331_n
  );


  buf

  (
    g1331_p_spl_,
    g1331_p
  );


  buf

  (
    g1330_n_spl_,
    g1330_n
  );


  buf

  (
    g1333_p_spl_,
    g1333_p
  );


  buf

  (
    g1330_p_spl_,
    g1330_p
  );


  buf

  (
    g1333_n_spl_,
    g1333_n
  );


  buf

  (
    lo038_buf_o2_p_spl_,
    lo038_buf_o2_p
  );


  buf

  (
    lo038_buf_o2_p_spl_0,
    lo038_buf_o2_p_spl_
  );


  buf

  (
    lo038_buf_o2_p_spl_00,
    lo038_buf_o2_p_spl_0
  );


  buf

  (
    lo038_buf_o2_p_spl_1,
    lo038_buf_o2_p_spl_
  );


  buf

  (
    lo038_buf_o2_n_spl_,
    lo038_buf_o2_n
  );


  buf

  (
    lo038_buf_o2_n_spl_0,
    lo038_buf_o2_n_spl_
  );


  buf

  (
    lo038_buf_o2_n_spl_1,
    lo038_buf_o2_n_spl_
  );


  buf

  (
    g1334_n_spl_,
    g1334_n
  );


  buf

  (
    g1334_p_spl_,
    g1334_p
  );


  buf

  (
    g1335_n_spl_,
    g1335_n
  );


  buf

  (
    g1337_p_spl_,
    g1337_p
  );


  buf

  (
    g1335_p_spl_,
    g1335_p
  );


  buf

  (
    g1337_n_spl_,
    g1337_n
  );


  buf

  (
    g1338_n_spl_,
    g1338_n
  );


  buf

  (
    g1338_p_spl_,
    g1338_p
  );


  buf

  (
    lo042_buf_o2_p_spl_,
    lo042_buf_o2_p
  );


  buf

  (
    lo042_buf_o2_p_spl_0,
    lo042_buf_o2_p_spl_
  );


  buf

  (
    lo042_buf_o2_p_spl_1,
    lo042_buf_o2_p_spl_
  );


  buf

  (
    lo042_buf_o2_n_spl_,
    lo042_buf_o2_n
  );


  buf

  (
    lo042_buf_o2_n_spl_0,
    lo042_buf_o2_n_spl_
  );


  buf

  (
    lo042_buf_o2_n_spl_1,
    lo042_buf_o2_n_spl_
  );


  buf

  (
    n1257_o2_n_spl_,
    n1257_o2_n
  );


  buf

  (
    n1281_o2_p_spl_,
    n1281_o2_p
  );


  buf

  (
    n1257_o2_p_spl_,
    n1257_o2_p
  );


  buf

  (
    n1281_o2_n_spl_,
    n1281_o2_n
  );


  buf

  (
    g1342_n_spl_,
    g1342_n
  );


  buf

  (
    g1342_p_spl_,
    g1342_p
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1345_n_spl_,
    g1345_n
  );


  buf

  (
    g1345_p_spl_,
    g1345_p
  );


  buf

  (
    g1340_n_spl_,
    g1340_n
  );


  buf

  (
    g1347_p_spl_,
    g1347_p
  );


  buf

  (
    g1340_p_spl_,
    g1340_p
  );


  buf

  (
    g1347_n_spl_,
    g1347_n
  );


  buf

  (
    g1348_n_spl_,
    g1348_n
  );


  buf

  (
    g1348_p_spl_,
    g1348_p
  );


  buf

  (
    g1339_n_spl_,
    g1339_n
  );


  buf

  (
    g1350_p_spl_,
    g1350_p
  );


  buf

  (
    g1339_p_spl_,
    g1339_p
  );


  buf

  (
    g1350_n_spl_,
    g1350_n
  );


  buf

  (
    g1351_n_spl_,
    g1351_n
  );


  buf

  (
    g1351_p_spl_,
    g1351_p
  );


  buf

  (
    g1352_n_spl_,
    g1352_n
  );


  buf

  (
    g1354_p_spl_,
    g1354_p
  );


  buf

  (
    g1352_p_spl_,
    g1352_p
  );


  buf

  (
    g1354_n_spl_,
    g1354_n
  );


  buf

  (
    g1355_n_spl_,
    g1355_n
  );


  buf

  (
    g1355_p_spl_,
    g1355_p
  );


  buf

  (
    lo046_buf_o2_p_spl_,
    lo046_buf_o2_p
  );


  buf

  (
    lo046_buf_o2_p_spl_0,
    lo046_buf_o2_p_spl_
  );


  buf

  (
    lo046_buf_o2_p_spl_1,
    lo046_buf_o2_p_spl_
  );


  buf

  (
    lo046_buf_o2_n_spl_,
    lo046_buf_o2_n
  );


  buf

  (
    lo046_buf_o2_n_spl_0,
    lo046_buf_o2_n_spl_
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1362_p_spl_,
    g1362_p
  );


  buf

  (
    g1360_p_spl_,
    g1360_p
  );


  buf

  (
    g1362_n_spl_,
    g1362_n
  );


  buf

  (
    g1363_n_spl_,
    g1363_n
  );


  buf

  (
    g1363_p_spl_,
    g1363_p
  );


  buf

  (
    g1359_n_spl_,
    g1359_n
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1359_p_spl_,
    g1359_p
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1366_n_spl_,
    g1366_n
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1358_n_spl_,
    g1358_n
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1358_p_spl_,
    g1358_p
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1369_n_spl_,
    g1369_n
  );


  buf

  (
    g1369_p_spl_,
    g1369_p
  );


  buf

  (
    g1357_n_spl_,
    g1357_n
  );


  buf

  (
    g1371_p_spl_,
    g1371_p
  );


  buf

  (
    g1357_p_spl_,
    g1357_p
  );


  buf

  (
    g1371_n_spl_,
    g1371_n
  );


  buf

  (
    g1372_n_spl_,
    g1372_n
  );


  buf

  (
    g1372_p_spl_,
    g1372_p
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1374_p_spl_,
    g1374_p
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1374_n_spl_,
    g1374_n
  );


  buf

  (
    g1375_n_spl_,
    g1375_n
  );


  buf

  (
    g1375_p_spl_,
    g1375_p
  );


  buf

  (
    g1376_n_spl_,
    g1376_n
  );


  buf

  (
    g1378_p_spl_,
    g1378_p
  );


  buf

  (
    g1376_p_spl_,
    g1376_p
  );


  buf

  (
    g1378_n_spl_,
    g1378_n
  );


  buf

  (
    g1379_n_spl_,
    g1379_n
  );


  buf

  (
    g1379_p_spl_,
    g1379_p
  );


  buf

  (
    g1384_n_spl_,
    g1384_n
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1384_p_spl_,
    g1384_p
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1387_n_spl_,
    g1387_n
  );


  buf

  (
    g1387_p_spl_,
    g1387_p
  );


  buf

  (
    g1383_n_spl_,
    g1383_n
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1383_p_spl_,
    g1383_p
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1390_n_spl_,
    g1390_n
  );


  buf

  (
    g1390_p_spl_,
    g1390_p
  );


  buf

  (
    g1382_n_spl_,
    g1382_n
  );


  buf

  (
    g1392_p_spl_,
    g1392_p
  );


  buf

  (
    g1382_p_spl_,
    g1382_p
  );


  buf

  (
    g1392_n_spl_,
    g1392_n
  );


  buf

  (
    g1393_n_spl_,
    g1393_n
  );


  buf

  (
    g1393_p_spl_,
    g1393_p
  );


  buf

  (
    g1381_n_spl_,
    g1381_n
  );


  buf

  (
    g1395_p_spl_,
    g1395_p
  );


  buf

  (
    g1381_p_spl_,
    g1381_p
  );


  buf

  (
    g1395_n_spl_,
    g1395_n
  );


  buf

  (
    g1396_n_spl_,
    g1396_n
  );


  buf

  (
    g1396_p_spl_,
    g1396_p
  );


  buf

  (
    g1380_n_spl_,
    g1380_n
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1380_p_spl_,
    g1380_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1250_p_spl_,
    g1250_p
  );


  buf

  (
    g1016_p_spl_,
    g1016_p
  );


  buf

  (
    n2833_lo_n_spl_,
    n2833_lo_n
  );


  buf

  (
    n2833_lo_n_spl_0,
    n2833_lo_n_spl_
  );


  buf

  (
    n2833_lo_n_spl_00,
    n2833_lo_n_spl_0
  );


  buf

  (
    n2833_lo_n_spl_1,
    n2833_lo_n_spl_
  );


  buf

  (
    n2770_lo_n_spl_,
    n2770_lo_n
  );


  buf

  (
    n2770_lo_n_spl_0,
    n2770_lo_n_spl_
  );


  buf

  (
    n2770_lo_n_spl_00,
    n2770_lo_n_spl_0
  );


  buf

  (
    n2770_lo_n_spl_000,
    n2770_lo_n_spl_00
  );


  buf

  (
    n2770_lo_n_spl_001,
    n2770_lo_n_spl_00
  );


  buf

  (
    n2770_lo_n_spl_01,
    n2770_lo_n_spl_0
  );


  buf

  (
    n2770_lo_n_spl_010,
    n2770_lo_n_spl_01
  );


  buf

  (
    n2770_lo_n_spl_1,
    n2770_lo_n_spl_
  );


  buf

  (
    n2770_lo_n_spl_10,
    n2770_lo_n_spl_1
  );


  buf

  (
    n2770_lo_n_spl_11,
    n2770_lo_n_spl_1
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_000,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_001,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_01,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_010,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_011,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_10,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_100,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_101,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_11,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_110,
    G20_n_spl_11
  );


  buf

  (
    g946_n_spl_,
    g946_n
  );


  buf

  (
    g1404_n_spl_,
    g1404_n
  );


  buf

  (
    g1406_p_spl_,
    g1406_p
  );


  buf

  (
    g934_n_spl_,
    g934_n
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1411_p_spl_,
    g1411_p
  );


  buf

  (
    g922_n_spl_,
    g922_n
  );


  buf

  (
    g1414_n_spl_,
    g1414_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g1419_n_spl_,
    g1419_n
  );


  buf

  (
    g1421_p_spl_,
    g1421_p
  );


  buf

  (
    g915_n_spl_,
    g915_n
  );


  buf

  (
    g1424_n_spl_,
    g1424_n
  );


  buf

  (
    g1426_p_spl_,
    g1426_p
  );


  buf

  (
    g911_n_spl_,
    g911_n
  );


  buf

  (
    g1429_n_spl_,
    g1429_n
  );


  buf

  (
    g1431_p_spl_,
    g1431_p
  );


  buf

  (
    g1013_n_spl_,
    g1013_n
  );


  buf

  (
    g1015_p_spl_,
    g1015_p
  );


  buf

  (
    n2833_lo_p_spl_,
    n2833_lo_p
  );


  buf

  (
    n2833_lo_p_spl_0,
    n2833_lo_p_spl_
  );


  buf

  (
    n2833_lo_p_spl_00,
    n2833_lo_p_spl_0
  );


  buf

  (
    n2833_lo_p_spl_1,
    n2833_lo_p_spl_
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1107_n_spl_,
    g1107_n
  );


  buf

  (
    g1053_n_spl_,
    g1053_n
  );


  buf

  (
    g1459_n_spl_,
    g1459_n
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1459_p_spl_,
    g1459_p
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1462_n_spl_,
    g1462_n
  );


  buf

  (
    g1462_p_spl_,
    g1462_p
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1464_n_spl_,
    g1464_n
  );


  buf

  (
    g1465_n_spl_,
    g1465_n
  );


  buf

  (
    g1465_p_spl_,
    g1465_p
  );


  buf

  (
    g1457_n_spl_,
    g1457_n
  );


  buf

  (
    g1467_p_spl_,
    g1467_p
  );


  buf

  (
    g1457_p_spl_,
    g1457_p
  );


  buf

  (
    g1467_n_spl_,
    g1467_n
  );


  buf

  (
    g1468_n_spl_,
    g1468_n
  );


  buf

  (
    g1468_p_spl_,
    g1468_p
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1456_p_spl_,
    g1456_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1455_n_spl_,
    g1455_n
  );


  buf

  (
    g1473_p_spl_,
    g1473_p
  );


  buf

  (
    g1454_n_spl_,
    g1454_n
  );


  buf

  (
    g1476_p_spl_,
    g1476_p
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1482_p_spl_,
    g1482_p
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1479_n_spl_,
    g1479_n
  );


  buf

  (
    g1485_p_spl_,
    g1485_p
  );


  buf

  (
    g1479_p_spl_,
    g1479_p
  );


  buf

  (
    g1485_n_spl_,
    g1485_n
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1492_n_spl_,
    g1492_n
  );


  buf

  (
    g1494_p_spl_,
    g1494_p
  );


  buf

  (
    g1492_p_spl_,
    g1492_p
  );


  buf

  (
    g1494_n_spl_,
    g1494_n
  );


  buf

  (
    g1495_n_spl_,
    g1495_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1497_p_spl_,
    g1497_p
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1497_n_spl_,
    g1497_n
  );


  buf

  (
    g1498_n_spl_,
    g1498_n
  );


  buf

  (
    g1504_n_spl_,
    g1504_n
  );


  buf

  (
    g1506_p_spl_,
    g1506_p
  );


  buf

  (
    g1504_p_spl_,
    g1504_p
  );


  buf

  (
    g1506_n_spl_,
    g1506_n
  );


  buf

  (
    g1507_n_spl_,
    g1507_n
  );


  buf

  (
    g1503_n_spl_,
    g1503_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1503_p_spl_,
    g1503_p
  );


  buf

  (
    g1509_n_spl_,
    g1509_n
  );


  buf

  (
    g1510_n_spl_,
    g1510_n
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    n2770_lo_p_spl_,
    n2770_lo_p
  );


  buf

  (
    n2770_lo_p_spl_0,
    n2770_lo_p_spl_
  );


  buf

  (
    n2770_lo_p_spl_00,
    n2770_lo_p_spl_0
  );


  buf

  (
    n2770_lo_p_spl_000,
    n2770_lo_p_spl_00
  );


  buf

  (
    n2770_lo_p_spl_001,
    n2770_lo_p_spl_00
  );


  buf

  (
    n2770_lo_p_spl_01,
    n2770_lo_p_spl_0
  );


  buf

  (
    n2770_lo_p_spl_1,
    n2770_lo_p_spl_
  );


  buf

  (
    n2770_lo_p_spl_10,
    n2770_lo_p_spl_1
  );


  buf

  (
    n2770_lo_p_spl_11,
    n2770_lo_p_spl_1
  );


  buf

  (
    g1399_n_spl_,
    g1399_n
  );


  buf

  (
    g1328_n_spl_,
    g1328_n
  );


  buf

  (
    g1526_n_spl_,
    g1526_n
  );


  buf

  (
    g1527_n_spl_,
    g1527_n
  );


  buf

  (
    g1526_p_spl_,
    g1526_p
  );


  buf

  (
    g1527_p_spl_,
    g1527_p
  );


  buf

  (
    g1528_p_spl_,
    g1528_p
  );


  buf

  (
    g1525_n_spl_,
    g1525_n
  );


  buf

  (
    g1530_p_spl_,
    g1530_p
  );


  buf

  (
    g1525_p_spl_,
    g1525_p
  );


  buf

  (
    g1530_n_spl_,
    g1530_n
  );


  buf

  (
    g1531_p_spl_,
    g1531_p
  );


  buf

  (
    g1537_n_spl_,
    g1537_n
  );


  buf

  (
    g1539_p_spl_,
    g1539_p
  );


  buf

  (
    g1537_p_spl_,
    g1537_p
  );


  buf

  (
    g1539_n_spl_,
    g1539_n
  );


  buf

  (
    g1540_p_spl_,
    g1540_p
  );


  buf

  (
    g1536_n_spl_,
    g1536_n
  );


  buf

  (
    g1542_p_spl_,
    g1542_p
  );


  buf

  (
    g1536_p_spl_,
    g1536_p
  );


  buf

  (
    g1542_n_spl_,
    g1542_n
  );


  buf

  (
    g1543_p_spl_,
    g1543_p
  );


  buf

  (
    g1242_p_spl_,
    g1242_p
  );


  buf

  (
    lo014_buf_o2_p_spl_,
    lo014_buf_o2_p
  );


  buf

  (
    lo014_buf_o2_p_spl_0,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_p_spl_00,
    lo014_buf_o2_p_spl_0
  );


  buf

  (
    lo014_buf_o2_p_spl_1,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_n_spl_,
    lo014_buf_o2_n
  );


  buf

  (
    lo014_buf_o2_n_spl_0,
    lo014_buf_o2_n_spl_
  );


  buf

  (
    lo014_buf_o2_n_spl_1,
    lo014_buf_o2_n_spl_
  );


  buf

  (
    n655_o2_n_spl_,
    n655_o2_n
  );


  buf

  (
    n679_o2_p_spl_,
    n679_o2_p
  );


  buf

  (
    n655_o2_p_spl_,
    n655_o2_p
  );


  buf

  (
    n679_o2_n_spl_,
    n679_o2_n
  );


  buf

  (
    g1554_n_spl_,
    g1554_n
  );


  buf

  (
    g1554_p_spl_,
    g1554_p
  );


  buf

  (
    g1553_n_spl_,
    g1553_n
  );


  buf

  (
    g1556_p_spl_,
    g1556_p
  );


  buf

  (
    g1553_p_spl_,
    g1553_p
  );


  buf

  (
    g1556_n_spl_,
    g1556_n
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    g1557_p_spl_,
    g1557_p
  );


  buf

  (
    g1552_n_spl_,
    g1552_n
  );


  buf

  (
    g1559_p_spl_,
    g1559_p
  );


  buf

  (
    g1552_p_spl_,
    g1552_p
  );


  buf

  (
    g1559_n_spl_,
    g1559_n
  );


  buf

  (
    g1560_n_spl_,
    g1560_n
  );


  buf

  (
    g1560_p_spl_,
    g1560_p
  );


  buf

  (
    g1551_n_spl_,
    g1551_n
  );


  buf

  (
    g1562_p_spl_,
    g1562_p
  );


  buf

  (
    g1551_p_spl_,
    g1551_p
  );


  buf

  (
    g1562_n_spl_,
    g1562_n
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1563_p_spl_,
    g1563_p
  );


  buf

  (
    g1550_n_spl_,
    g1550_n
  );


  buf

  (
    g1565_p_spl_,
    g1565_p
  );


  buf

  (
    g1550_p_spl_,
    g1550_p
  );


  buf

  (
    g1565_n_spl_,
    g1565_n
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1566_p_spl_,
    g1566_p
  );


  buf

  (
    g1549_n_spl_,
    g1549_n
  );


  buf

  (
    g1568_p_spl_,
    g1568_p
  );


  buf

  (
    g1549_p_spl_,
    g1549_p
  );


  buf

  (
    g1568_n_spl_,
    g1568_n
  );


  buf

  (
    g1569_n_spl_,
    g1569_n
  );


  buf

  (
    g1569_p_spl_,
    g1569_p
  );


  buf

  (
    g1548_n_spl_,
    g1548_n
  );


  buf

  (
    g1571_p_spl_,
    g1571_p
  );


  buf

  (
    g1548_p_spl_,
    g1548_p
  );


  buf

  (
    g1571_n_spl_,
    g1571_n
  );


  buf

  (
    g1572_n_spl_,
    g1572_n
  );


  buf

  (
    g1572_p_spl_,
    g1572_p
  );


  buf

  (
    g1547_n_spl_,
    g1547_n
  );


  buf

  (
    g1574_p_spl_,
    g1574_p
  );


  buf

  (
    g1400_p_spl_,
    g1400_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    g1580_p_spl_,
    g1580_p
  );


  buf

  (
    g1581_p_spl_,
    g1581_p
  );


  buf

  (
    g1580_n_spl_,
    g1580_n
  );


  buf

  (
    g1581_n_spl_,
    g1581_n
  );


  buf

  (
    g1582_n_spl_,
    g1582_n
  );


  buf

  (
    g1582_n_spl_0,
    g1582_n_spl_
  );


  buf

  (
    g1582_p_spl_,
    g1582_p
  );


  buf

  (
    g1582_p_spl_0,
    g1582_p_spl_
  );


  buf

  (
    g1584_n_spl_,
    g1584_n
  );


  buf

  (
    g1584_p_spl_,
    g1584_p
  );


  buf

  (
    g1585_n_spl_,
    g1585_n
  );


  buf

  (
    g1585_p_spl_,
    g1585_p
  );


  buf

  (
    g1579_n_spl_,
    g1579_n
  );


  buf

  (
    g1587_p_spl_,
    g1587_p
  );


  buf

  (
    g1579_p_spl_,
    g1579_p
  );


  buf

  (
    g1587_n_spl_,
    g1587_n
  );


  buf

  (
    g1588_n_spl_,
    g1588_n
  );


  buf

  (
    g1588_p_spl_,
    g1588_p
  );


  buf

  (
    g1578_n_spl_,
    g1578_n
  );


  buf

  (
    g1590_p_spl_,
    g1590_p
  );


  buf

  (
    g1603_n_spl_,
    g1603_n
  );


  buf

  (
    g1605_p_spl_,
    g1605_p
  );


  buf

  (
    g1603_p_spl_,
    g1603_p
  );


  buf

  (
    g1605_n_spl_,
    g1605_n
  );


  buf

  (
    g1606_n_spl_,
    g1606_n
  );


  buf

  (
    g1606_p_spl_,
    g1606_p
  );


  buf

  (
    g1602_n_spl_,
    g1602_n
  );


  buf

  (
    g1608_p_spl_,
    g1608_p
  );


  buf

  (
    g1602_p_spl_,
    g1602_p
  );


  buf

  (
    g1608_n_spl_,
    g1608_n
  );


  buf

  (
    g1609_n_spl_,
    g1609_n
  );


  buf

  (
    g1609_p_spl_,
    g1609_p
  );


  buf

  (
    g1601_n_spl_,
    g1601_n
  );


  buf

  (
    g1611_p_spl_,
    g1611_p
  );


  buf

  (
    g1601_p_spl_,
    g1601_p
  );


  buf

  (
    g1611_n_spl_,
    g1611_n
  );


  buf

  (
    g1612_n_spl_,
    g1612_n
  );


  buf

  (
    g1616_n_spl_,
    g1616_n
  );


  buf

  (
    g1618_n_spl_,
    g1618_n
  );


  buf

  (
    g1620_p_spl_,
    g1620_p
  );


  buf

  (
    g1618_p_spl_,
    g1618_p
  );


  buf

  (
    g1620_n_spl_,
    g1620_n
  );


  buf

  (
    g1621_n_spl_,
    g1621_n
  );


  buf

  (
    g1625_n_spl_,
    g1625_n
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1515_p_spl_,
    g1515_p
  );


  buf

  (
    g1402_n_spl_,
    g1402_n
  );


  buf

  (
    g1577_p_spl_,
    g1577_p
  );


  buf

  (
    g1403_n_spl_,
    g1403_n
  );


  buf

  (
    g1593_p_spl_,
    g1593_p
  );


  buf

  (
    g1438_n_spl_,
    g1438_n
  );


  buf

  (
    g1442_n_spl_,
    g1442_n
  );


  buf

  (
    g1446_n_spl_,
    g1446_n
  );


  buf

  (
    g1450_n_spl_,
    g1450_n
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1489_n_spl_,
    g1489_n
  );


  buf

  (
    g1501_n_spl_,
    g1501_n
  );


  buf

  (
    g1513_n_spl_,
    g1513_n
  );


  buf

  (
    g1630_p_spl_,
    g1630_p
  );


  buf

  (
    lo018_buf_o2_p_spl_,
    lo018_buf_o2_p
  );


  buf

  (
    lo018_buf_o2_p_spl_0,
    lo018_buf_o2_p_spl_
  );


  buf

  (
    lo018_buf_o2_p_spl_00,
    lo018_buf_o2_p_spl_0
  );


  buf

  (
    lo018_buf_o2_p_spl_1,
    lo018_buf_o2_p_spl_
  );


  buf

  (
    lo018_buf_o2_n_spl_,
    lo018_buf_o2_n
  );


  buf

  (
    lo018_buf_o2_n_spl_0,
    lo018_buf_o2_n_spl_
  );


  buf

  (
    lo018_buf_o2_n_spl_1,
    lo018_buf_o2_n_spl_
  );


  buf

  (
    n717_o2_n_spl_,
    n717_o2_n
  );


  buf

  (
    n741_o2_p_spl_,
    n741_o2_p
  );


  buf

  (
    n717_o2_p_spl_,
    n717_o2_p
  );


  buf

  (
    n741_o2_n_spl_,
    n741_o2_n
  );


  buf

  (
    g1661_n_spl_,
    g1661_n
  );


  buf

  (
    g1661_p_spl_,
    g1661_p
  );


  buf

  (
    g1660_n_spl_,
    g1660_n
  );


  buf

  (
    g1663_p_spl_,
    g1663_p
  );


  buf

  (
    g1660_p_spl_,
    g1660_p
  );


  buf

  (
    g1663_n_spl_,
    g1663_n
  );


  buf

  (
    g1664_n_spl_,
    g1664_n
  );


  buf

  (
    g1664_p_spl_,
    g1664_p
  );


  buf

  (
    g1659_n_spl_,
    g1659_n
  );


  buf

  (
    g1666_p_spl_,
    g1666_p
  );


  buf

  (
    g1659_p_spl_,
    g1659_p
  );


  buf

  (
    g1666_n_spl_,
    g1666_n
  );


  buf

  (
    g1667_n_spl_,
    g1667_n
  );


  buf

  (
    g1667_p_spl_,
    g1667_p
  );


  buf

  (
    g1658_n_spl_,
    g1658_n
  );


  buf

  (
    g1669_p_spl_,
    g1669_p
  );


  buf

  (
    g1658_p_spl_,
    g1658_p
  );


  buf

  (
    g1669_n_spl_,
    g1669_n
  );


  buf

  (
    g1670_n_spl_,
    g1670_n
  );


  buf

  (
    g1670_p_spl_,
    g1670_p
  );


  buf

  (
    g1657_n_spl_,
    g1657_n
  );


  buf

  (
    g1672_p_spl_,
    g1672_p
  );


  buf

  (
    g1657_p_spl_,
    g1657_p
  );


  buf

  (
    g1672_n_spl_,
    g1672_n
  );


  buf

  (
    g1673_n_spl_,
    g1673_n
  );


  buf

  (
    g1673_p_spl_,
    g1673_p
  );


  buf

  (
    g1656_n_spl_,
    g1656_n
  );


  buf

  (
    g1675_p_spl_,
    g1675_p
  );


  buf

  (
    g1656_p_spl_,
    g1656_p
  );


  buf

  (
    g1675_n_spl_,
    g1675_n
  );


  buf

  (
    g1676_n_spl_,
    g1676_n
  );


  buf

  (
    g1676_p_spl_,
    g1676_p
  );


  buf

  (
    g1655_n_spl_,
    g1655_n
  );


  buf

  (
    g1678_p_spl_,
    g1678_p
  );


  buf

  (
    g1655_p_spl_,
    g1655_p
  );


  buf

  (
    g1678_n_spl_,
    g1678_n
  );


  buf

  (
    g1679_n_spl_,
    g1679_n
  );


  buf

  (
    g1679_p_spl_,
    g1679_p
  );


  buf

  (
    g1654_n_spl_,
    g1654_n
  );


  buf

  (
    g1681_p_spl_,
    g1681_p
  );


  buf

  (
    g1654_p_spl_,
    g1654_p
  );


  buf

  (
    g1681_n_spl_,
    g1681_n
  );


  buf

  (
    g1682_n_spl_,
    g1682_n
  );


  buf

  (
    g1685_n_spl_,
    g1685_n
  );


  buf

  (
    g1546_n_spl_,
    g1546_n
  );


  buf

  (
    g1688_n_spl_,
    g1688_n
  );


  buf

  (
    g1690_p_spl_,
    g1690_p
  );


  buf

  (
    g1534_n_spl_,
    g1534_n
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1695_p_spl_,
    g1695_p
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1523_n_spl_,
    g1523_n
  );


  buf

  (
    g1702_n_spl_,
    g1702_n
  );


  buf

  (
    g1704_p_spl_,
    g1704_p
  );


  buf

  (
    lo022_buf_o2_p_spl_,
    lo022_buf_o2_p
  );


  buf

  (
    lo022_buf_o2_p_spl_0,
    lo022_buf_o2_p_spl_
  );


  buf

  (
    lo022_buf_o2_p_spl_00,
    lo022_buf_o2_p_spl_0
  );


  buf

  (
    lo022_buf_o2_p_spl_1,
    lo022_buf_o2_p_spl_
  );


  buf

  (
    lo022_buf_o2_n_spl_,
    lo022_buf_o2_n
  );


  buf

  (
    lo022_buf_o2_n_spl_0,
    lo022_buf_o2_n_spl_
  );


  buf

  (
    lo022_buf_o2_n_spl_1,
    lo022_buf_o2_n_spl_
  );


  buf

  (
    n787_o2_n_spl_,
    n787_o2_n
  );


  buf

  (
    n811_o2_p_spl_,
    n811_o2_p
  );


  buf

  (
    n787_o2_p_spl_,
    n787_o2_p
  );


  buf

  (
    n811_o2_n_spl_,
    n811_o2_n
  );


  buf

  (
    g1714_n_spl_,
    g1714_n
  );


  buf

  (
    g1714_p_spl_,
    g1714_p
  );


  buf

  (
    g1713_n_spl_,
    g1713_n
  );


  buf

  (
    g1716_p_spl_,
    g1716_p
  );


  buf

  (
    g1713_p_spl_,
    g1713_p
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1717_n_spl_,
    g1717_n
  );


  buf

  (
    g1717_p_spl_,
    g1717_p
  );


  buf

  (
    g1712_n_spl_,
    g1712_n
  );


  buf

  (
    g1719_p_spl_,
    g1719_p
  );


  buf

  (
    g1712_p_spl_,
    g1712_p
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


  buf

  (
    g1720_n_spl_,
    g1720_n
  );


  buf

  (
    g1720_p_spl_,
    g1720_p
  );


  buf

  (
    g1711_n_spl_,
    g1711_n
  );


  buf

  (
    g1722_p_spl_,
    g1722_p
  );


  buf

  (
    g1711_p_spl_,
    g1711_p
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1723_n_spl_,
    g1723_n
  );


  buf

  (
    g1723_p_spl_,
    g1723_p
  );


  buf

  (
    g1710_n_spl_,
    g1710_n
  );


  buf

  (
    g1725_p_spl_,
    g1725_p
  );


  buf

  (
    g1710_p_spl_,
    g1710_p
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1726_n_spl_,
    g1726_n
  );


  buf

  (
    g1726_p_spl_,
    g1726_p
  );


  buf

  (
    g1709_n_spl_,
    g1709_n
  );


  buf

  (
    g1728_p_spl_,
    g1728_p
  );


  buf

  (
    g1709_p_spl_,
    g1709_p
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    g1729_n_spl_,
    g1729_n
  );


  buf

  (
    g1729_p_spl_,
    g1729_p
  );


  buf

  (
    g1708_n_spl_,
    g1708_n
  );


  buf

  (
    g1731_p_spl_,
    g1731_p
  );


  buf

  (
    g1708_p_spl_,
    g1708_p
  );


  buf

  (
    g1731_n_spl_,
    g1731_n
  );


  buf

  (
    g1732_n_spl_,
    g1732_n
  );


  buf

  (
    g1732_p_spl_,
    g1732_p
  );


  buf

  (
    g1707_n_spl_,
    g1707_n
  );


  buf

  (
    g1734_p_spl_,
    g1734_p
  );


  buf

  (
    g1707_p_spl_,
    g1707_p
  );


  buf

  (
    g1734_n_spl_,
    g1734_n
  );


  buf

  (
    g1735_p_spl_,
    g1735_p
  );


  buf

  (
    g1739_p_spl_,
    g1739_p
  );


  buf

  (
    lo026_buf_o2_p_spl_,
    lo026_buf_o2_p
  );


  buf

  (
    lo026_buf_o2_p_spl_0,
    lo026_buf_o2_p_spl_
  );


  buf

  (
    lo026_buf_o2_p_spl_00,
    lo026_buf_o2_p_spl_0
  );


  buf

  (
    lo026_buf_o2_p_spl_1,
    lo026_buf_o2_p_spl_
  );


  buf

  (
    lo026_buf_o2_n_spl_,
    lo026_buf_o2_n
  );


  buf

  (
    lo026_buf_o2_n_spl_0,
    lo026_buf_o2_n_spl_
  );


  buf

  (
    lo026_buf_o2_n_spl_1,
    lo026_buf_o2_n_spl_
  );


  buf

  (
    n865_o2_n_spl_,
    n865_o2_n
  );


  buf

  (
    n889_o2_p_spl_,
    n889_o2_p
  );


  buf

  (
    n865_o2_p_spl_,
    n865_o2_p
  );


  buf

  (
    n889_o2_n_spl_,
    n889_o2_n
  );


  buf

  (
    g1749_n_spl_,
    g1749_n
  );


  buf

  (
    g1749_p_spl_,
    g1749_p
  );


  buf

  (
    g1748_n_spl_,
    g1748_n
  );


  buf

  (
    g1751_p_spl_,
    g1751_p
  );


  buf

  (
    g1748_p_spl_,
    g1748_p
  );


  buf

  (
    g1751_n_spl_,
    g1751_n
  );


  buf

  (
    g1752_n_spl_,
    g1752_n
  );


  buf

  (
    g1752_p_spl_,
    g1752_p
  );


  buf

  (
    g1747_n_spl_,
    g1747_n
  );


  buf

  (
    g1754_p_spl_,
    g1754_p
  );


  buf

  (
    g1747_p_spl_,
    g1747_p
  );


  buf

  (
    g1754_n_spl_,
    g1754_n
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1755_p_spl_,
    g1755_p
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1757_p_spl_,
    g1757_p
  );


  buf

  (
    g1746_p_spl_,
    g1746_p
  );


  buf

  (
    g1757_n_spl_,
    g1757_n
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1745_n_spl_,
    g1745_n
  );


  buf

  (
    g1760_p_spl_,
    g1760_p
  );


  buf

  (
    g1745_p_spl_,
    g1745_p
  );


  buf

  (
    g1760_n_spl_,
    g1760_n
  );


  buf

  (
    g1761_n_spl_,
    g1761_n
  );


  buf

  (
    g1761_p_spl_,
    g1761_p
  );


  buf

  (
    g1744_n_spl_,
    g1744_n
  );


  buf

  (
    g1763_p_spl_,
    g1763_p
  );


  buf

  (
    g1744_p_spl_,
    g1744_p
  );


  buf

  (
    g1763_n_spl_,
    g1763_n
  );


  buf

  (
    g1764_n_spl_,
    g1764_n
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1743_n_spl_,
    g1743_n
  );


  buf

  (
    g1766_p_spl_,
    g1766_p
  );


  buf

  (
    g1743_p_spl_,
    g1743_p
  );


  buf

  (
    g1766_n_spl_,
    g1766_n
  );


  buf

  (
    g1767_n_spl_,
    g1767_n
  );


  buf

  (
    g1767_p_spl_,
    g1767_p
  );


  buf

  (
    g1742_n_spl_,
    g1742_n
  );


  buf

  (
    g1769_p_spl_,
    g1769_p
  );


  buf

  (
    g1742_p_spl_,
    g1742_p
  );


  buf

  (
    g1769_n_spl_,
    g1769_n
  );


  buf

  (
    g1770_p_spl_,
    g1770_p
  );


  buf

  (
    g1741_n_spl_,
    g1741_n
  );


  buf

  (
    g1772_p_spl_,
    g1772_p
  );


  buf

  (
    g1740_n_spl_,
    g1740_n
  );


  buf

  (
    g1775_p_spl_,
    g1775_p
  );


  buf

  (
    lo030_buf_o2_p_spl_,
    lo030_buf_o2_p
  );


  buf

  (
    lo030_buf_o2_p_spl_0,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    lo030_buf_o2_p_spl_00,
    lo030_buf_o2_p_spl_0
  );


  buf

  (
    lo030_buf_o2_p_spl_1,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    lo030_buf_o2_n_spl_,
    lo030_buf_o2_n
  );


  buf

  (
    lo030_buf_o2_n_spl_0,
    lo030_buf_o2_n_spl_
  );


  buf

  (
    lo030_buf_o2_n_spl_1,
    lo030_buf_o2_n_spl_
  );


  buf

  (
    n951_o2_n_spl_,
    n951_o2_n
  );


  buf

  (
    n975_o2_p_spl_,
    n975_o2_p
  );


  buf

  (
    n951_o2_p_spl_,
    n951_o2_p
  );


  buf

  (
    n975_o2_n_spl_,
    n975_o2_n
  );


  buf

  (
    g1787_n_spl_,
    g1787_n
  );


  buf

  (
    g1787_p_spl_,
    g1787_p
  );


  buf

  (
    g1786_n_spl_,
    g1786_n
  );


  buf

  (
    g1789_p_spl_,
    g1789_p
  );


  buf

  (
    g1786_p_spl_,
    g1786_p
  );


  buf

  (
    g1789_n_spl_,
    g1789_n
  );


  buf

  (
    g1790_n_spl_,
    g1790_n
  );


  buf

  (
    g1790_p_spl_,
    g1790_p
  );


  buf

  (
    g1785_n_spl_,
    g1785_n
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    g1792_n_spl_,
    g1792_n
  );


  buf

  (
    g1793_n_spl_,
    g1793_n
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1784_n_spl_,
    g1784_n
  );


  buf

  (
    g1795_p_spl_,
    g1795_p
  );


  buf

  (
    g1784_p_spl_,
    g1784_p
  );


  buf

  (
    g1795_n_spl_,
    g1795_n
  );


  buf

  (
    g1796_n_spl_,
    g1796_n
  );


  buf

  (
    g1796_p_spl_,
    g1796_p
  );


  buf

  (
    g1783_n_spl_,
    g1783_n
  );


  buf

  (
    g1798_p_spl_,
    g1798_p
  );


  buf

  (
    g1783_p_spl_,
    g1783_p
  );


  buf

  (
    g1798_n_spl_,
    g1798_n
  );


  buf

  (
    g1799_n_spl_,
    g1799_n
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1782_n_spl_,
    g1782_n
  );


  buf

  (
    g1801_p_spl_,
    g1801_p
  );


  buf

  (
    g1782_p_spl_,
    g1782_p
  );


  buf

  (
    g1801_n_spl_,
    g1801_n
  );


  buf

  (
    g1802_n_spl_,
    g1802_n
  );


  buf

  (
    g1802_p_spl_,
    g1802_p
  );


  buf

  (
    g1781_n_spl_,
    g1781_n
  );


  buf

  (
    g1804_p_spl_,
    g1804_p
  );


  buf

  (
    g1781_p_spl_,
    g1781_p
  );


  buf

  (
    g1804_n_spl_,
    g1804_n
  );


  buf

  (
    g1805_n_spl_,
    g1805_n
  );


  buf

  (
    g1805_p_spl_,
    g1805_p
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1807_p_spl_,
    g1807_p
  );


  buf

  (
    g1780_p_spl_,
    g1780_p
  );


  buf

  (
    g1807_n_spl_,
    g1807_n
  );


  buf

  (
    g1808_p_spl_,
    g1808_p
  );


  buf

  (
    g1779_n_spl_,
    g1779_n
  );


  buf

  (
    g1810_p_spl_,
    g1810_p
  );


  buf

  (
    g1778_n_spl_,
    g1778_n
  );


  buf

  (
    g1813_p_spl_,
    g1813_p
  );


  buf

  (
    lo034_buf_o2_p_spl_,
    lo034_buf_o2_p
  );


  buf

  (
    lo034_buf_o2_p_spl_0,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    lo034_buf_o2_p_spl_00,
    lo034_buf_o2_p_spl_0
  );


  buf

  (
    lo034_buf_o2_p_spl_1,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    lo034_buf_o2_n_spl_,
    lo034_buf_o2_n
  );


  buf

  (
    lo034_buf_o2_n_spl_0,
    lo034_buf_o2_n_spl_
  );


  buf

  (
    lo034_buf_o2_n_spl_1,
    lo034_buf_o2_n_spl_
  );


  buf

  (
    g1824_n_spl_,
    g1824_n
  );


  buf

  (
    g1826_p_spl_,
    g1826_p
  );


  buf

  (
    g1824_p_spl_,
    g1824_p
  );


  buf

  (
    g1826_n_spl_,
    g1826_n
  );


  buf

  (
    g1827_n_spl_,
    g1827_n
  );


  buf

  (
    g1827_p_spl_,
    g1827_p
  );


  buf

  (
    g1823_n_spl_,
    g1823_n
  );


  buf

  (
    g1829_p_spl_,
    g1829_p
  );


  buf

  (
    g1823_p_spl_,
    g1823_p
  );


  buf

  (
    g1829_n_spl_,
    g1829_n
  );


  buf

  (
    g1830_n_spl_,
    g1830_n
  );


  buf

  (
    g1830_p_spl_,
    g1830_p
  );


  buf

  (
    g1822_n_spl_,
    g1822_n
  );


  buf

  (
    g1832_p_spl_,
    g1832_p
  );


  buf

  (
    g1822_p_spl_,
    g1822_p
  );


  buf

  (
    g1832_n_spl_,
    g1832_n
  );


  buf

  (
    g1833_n_spl_,
    g1833_n
  );


  buf

  (
    g1833_p_spl_,
    g1833_p
  );


  buf

  (
    g1821_n_spl_,
    g1821_n
  );


  buf

  (
    g1835_p_spl_,
    g1835_p
  );


  buf

  (
    g1821_p_spl_,
    g1821_p
  );


  buf

  (
    g1835_n_spl_,
    g1835_n
  );


  buf

  (
    g1836_n_spl_,
    g1836_n
  );


  buf

  (
    g1836_p_spl_,
    g1836_p
  );


  buf

  (
    g1820_n_spl_,
    g1820_n
  );


  buf

  (
    g1838_p_spl_,
    g1838_p
  );


  buf

  (
    g1820_p_spl_,
    g1820_p
  );


  buf

  (
    g1838_n_spl_,
    g1838_n
  );


  buf

  (
    g1839_n_spl_,
    g1839_n
  );


  buf

  (
    g1839_p_spl_,
    g1839_p
  );


  buf

  (
    g1819_n_spl_,
    g1819_n
  );


  buf

  (
    g1841_p_spl_,
    g1841_p
  );


  buf

  (
    g1819_p_spl_,
    g1819_p
  );


  buf

  (
    g1841_n_spl_,
    g1841_n
  );


  buf

  (
    g1842_n_spl_,
    g1842_n
  );


  buf

  (
    g1842_p_spl_,
    g1842_p
  );


  buf

  (
    g1818_n_spl_,
    g1818_n
  );


  buf

  (
    g1844_p_spl_,
    g1844_p
  );


  buf

  (
    g1818_p_spl_,
    g1818_p
  );


  buf

  (
    g1844_n_spl_,
    g1844_n
  );


  buf

  (
    g1845_p_spl_,
    g1845_p
  );


  buf

  (
    g1817_n_spl_,
    g1817_n
  );


  buf

  (
    g1847_p_spl_,
    g1847_p
  );


  buf

  (
    g1816_n_spl_,
    g1816_n
  );


  buf

  (
    g1850_p_spl_,
    g1850_p
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1861_p_spl_,
    g1861_p
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1861_n_spl_,
    g1861_n
  );


  buf

  (
    g1862_n_spl_,
    g1862_n
  );


  buf

  (
    g1862_p_spl_,
    g1862_p
  );


  buf

  (
    g1858_n_spl_,
    g1858_n
  );


  buf

  (
    g1864_p_spl_,
    g1864_p
  );


  buf

  (
    g1858_p_spl_,
    g1858_p
  );


  buf

  (
    g1864_n_spl_,
    g1864_n
  );


  buf

  (
    g1865_n_spl_,
    g1865_n
  );


  buf

  (
    g1865_p_spl_,
    g1865_p
  );


  buf

  (
    g1857_n_spl_,
    g1857_n
  );


  buf

  (
    g1867_p_spl_,
    g1867_p
  );


  buf

  (
    g1857_p_spl_,
    g1857_p
  );


  buf

  (
    g1867_n_spl_,
    g1867_n
  );


  buf

  (
    g1868_n_spl_,
    g1868_n
  );


  buf

  (
    g1868_p_spl_,
    g1868_p
  );


  buf

  (
    g1856_n_spl_,
    g1856_n
  );


  buf

  (
    g1870_p_spl_,
    g1870_p
  );


  buf

  (
    g1856_p_spl_,
    g1856_p
  );


  buf

  (
    g1870_n_spl_,
    g1870_n
  );


  buf

  (
    g1871_n_spl_,
    g1871_n
  );


  buf

  (
    g1871_p_spl_,
    g1871_p
  );


  buf

  (
    g1855_n_spl_,
    g1855_n
  );


  buf

  (
    g1873_p_spl_,
    g1873_p
  );


  buf

  (
    g1855_p_spl_,
    g1855_p
  );


  buf

  (
    g1873_n_spl_,
    g1873_n
  );


  buf

  (
    g1874_p_spl_,
    g1874_p
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1876_p_spl_,
    g1876_p
  );


  buf

  (
    g1853_n_spl_,
    g1853_n
  );


  buf

  (
    g1879_p_spl_,
    g1879_p
  );


  buf

  (
    g1886_n_spl_,
    g1886_n
  );


  buf

  (
    g1888_p_spl_,
    g1888_p
  );


  buf

  (
    g1886_p_spl_,
    g1886_p
  );


  buf

  (
    g1888_n_spl_,
    g1888_n
  );


  buf

  (
    g1889_n_spl_,
    g1889_n
  );


  buf

  (
    g1889_p_spl_,
    g1889_p
  );


  buf

  (
    g1885_n_spl_,
    g1885_n
  );


  buf

  (
    g1891_p_spl_,
    g1891_p
  );


  buf

  (
    g1885_p_spl_,
    g1885_p
  );


  buf

  (
    g1891_n_spl_,
    g1891_n
  );


  buf

  (
    g1892_n_spl_,
    g1892_n
  );


  buf

  (
    g1892_p_spl_,
    g1892_p
  );


  buf

  (
    g1884_n_spl_,
    g1884_n
  );


  buf

  (
    g1894_p_spl_,
    g1894_p
  );


  buf

  (
    g1884_p_spl_,
    g1884_p
  );


  buf

  (
    g1894_n_spl_,
    g1894_n
  );


  buf

  (
    g1895_p_spl_,
    g1895_p
  );


  buf

  (
    g1883_n_spl_,
    g1883_n
  );


  buf

  (
    g1897_p_spl_,
    g1897_p
  );


  buf

  (
    g1882_n_spl_,
    g1882_n
  );


  buf

  (
    g1900_p_spl_,
    g1900_p
  );


  buf

  (
    g1905_n_spl_,
    g1905_n
  );


  buf

  (
    g1907_p_spl_,
    g1907_p
  );


  buf

  (
    g1905_p_spl_,
    g1905_p
  );


  buf

  (
    g1907_n_spl_,
    g1907_n
  );


  buf

  (
    g1908_p_spl_,
    g1908_p
  );


  buf

  (
    g1904_n_spl_,
    g1904_n
  );


  buf

  (
    g1910_p_spl_,
    g1910_p
  );


  buf

  (
    g1903_n_spl_,
    g1903_n
  );


  buf

  (
    g1913_p_spl_,
    g1913_p
  );


  buf

  (
    g1519_n_spl_,
    g1519_n
  );


  buf

  (
    g1916_n_spl_,
    g1916_n
  );


  buf

  (
    g1918_p_spl_,
    g1918_p
  );


  buf

  (
    g1921_p_spl_,
    g1921_p
  );


  buf

  (
    g1923_n_spl_,
    g1923_n
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_01,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    g1926_p_spl_,
    g1926_p
  );


  buf

  (
    g1927_p_spl_,
    g1927_p
  );


  buf

  (
    g1926_n_spl_,
    g1926_n
  );


  buf

  (
    g1927_n_spl_,
    g1927_n
  );


  buf

  (
    g1928_n_spl_,
    g1928_n
  );


  buf

  (
    g1928_n_spl_0,
    g1928_n_spl_
  );


  buf

  (
    g1928_p_spl_,
    g1928_p
  );


  buf

  (
    g1928_p_spl_0,
    g1928_p_spl_
  );


  buf

  (
    g1930_n_spl_,
    g1930_n
  );


  buf

  (
    g1930_p_spl_,
    g1930_p
  );


  buf

  (
    g1931_n_spl_,
    g1931_n
  );


  buf

  (
    g1931_p_spl_,
    g1931_p
  );


  buf

  (
    g1932_n_spl_,
    g1932_n
  );


  buf

  (
    g1934_p_spl_,
    g1934_p
  );


  buf

  (
    g1932_p_spl_,
    g1932_p
  );


  buf

  (
    g1934_n_spl_,
    g1934_n
  );


  buf

  (
    g1935_n_spl_,
    g1935_n
  );


  buf

  (
    g1935_p_spl_,
    g1935_p
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_01,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    g1938_p_spl_,
    g1938_p
  );


  buf

  (
    g1939_p_spl_,
    g1939_p
  );


  buf

  (
    g1938_n_spl_,
    g1938_n
  );


  buf

  (
    g1939_n_spl_,
    g1939_n
  );


  buf

  (
    g1940_n_spl_,
    g1940_n
  );


  buf

  (
    g1940_n_spl_0,
    g1940_n_spl_
  );


  buf

  (
    g1940_p_spl_,
    g1940_p
  );


  buf

  (
    g1940_p_spl_0,
    g1940_p_spl_
  );


  buf

  (
    g1942_n_spl_,
    g1942_n
  );


  buf

  (
    g1942_p_spl_,
    g1942_p
  );


  buf

  (
    g1943_n_spl_,
    g1943_n
  );


  buf

  (
    g1943_p_spl_,
    g1943_p
  );


  buf

  (
    g1937_n_spl_,
    g1937_n
  );


  buf

  (
    g1945_p_spl_,
    g1945_p
  );


  buf

  (
    g1937_p_spl_,
    g1937_p
  );


  buf

  (
    g1945_n_spl_,
    g1945_n
  );


  buf

  (
    g1946_n_spl_,
    g1946_n
  );


  buf

  (
    g1946_p_spl_,
    g1946_p
  );


  buf

  (
    g1936_n_spl_,
    g1936_n
  );


  buf

  (
    g1948_p_spl_,
    g1948_p
  );


  buf

  (
    g1936_p_spl_,
    g1936_p
  );


  buf

  (
    g1948_n_spl_,
    g1948_n
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_000,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_001,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_01,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_010,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_011,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_10,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_100,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_101,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_11,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_110,
    G20_p_spl_11
  );


  buf

  (
    g1949_n_spl_,
    g1949_n
  );


  buf

  (
    g1949_p_spl_,
    g1949_p
  );


  buf

  (
    g1950_n_spl_,
    g1950_n
  );


  buf

  (
    g1952_p_spl_,
    g1952_p
  );


  buf

  (
    g1950_p_spl_,
    g1950_p
  );


  buf

  (
    g1952_n_spl_,
    g1952_n
  );


  buf

  (
    g1953_n_spl_,
    g1953_n
  );


  buf

  (
    g1953_p_spl_,
    g1953_p
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_01,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    g1958_p_spl_,
    g1958_p
  );


  buf

  (
    g1959_p_spl_,
    g1959_p
  );


  buf

  (
    g1958_n_spl_,
    g1958_n
  );


  buf

  (
    g1959_n_spl_,
    g1959_n
  );


  buf

  (
    g1960_n_spl_,
    g1960_n
  );


  buf

  (
    g1960_n_spl_0,
    g1960_n_spl_
  );


  buf

  (
    g1960_p_spl_,
    g1960_p
  );


  buf

  (
    g1960_p_spl_0,
    g1960_p_spl_
  );


  buf

  (
    g1962_n_spl_,
    g1962_n
  );


  buf

  (
    g1962_p_spl_,
    g1962_p
  );


  buf

  (
    g1963_n_spl_,
    g1963_n
  );


  buf

  (
    g1963_p_spl_,
    g1963_p
  );


  buf

  (
    g1957_n_spl_,
    g1957_n
  );


  buf

  (
    g1965_p_spl_,
    g1965_p
  );


  buf

  (
    g1957_p_spl_,
    g1957_p
  );


  buf

  (
    g1965_n_spl_,
    g1965_n
  );


  buf

  (
    g1966_n_spl_,
    g1966_n
  );


  buf

  (
    g1966_p_spl_,
    g1966_p
  );


  buf

  (
    g1956_n_spl_,
    g1956_n
  );


  buf

  (
    g1968_p_spl_,
    g1968_p
  );


  buf

  (
    g1956_p_spl_,
    g1956_p
  );


  buf

  (
    g1968_n_spl_,
    g1968_n
  );


  buf

  (
    g1969_n_spl_,
    g1969_n
  );


  buf

  (
    g1969_p_spl_,
    g1969_p
  );


  buf

  (
    g1955_n_spl_,
    g1955_n
  );


  buf

  (
    g1971_p_spl_,
    g1971_p
  );


  buf

  (
    g1955_p_spl_,
    g1955_p
  );


  buf

  (
    g1971_n_spl_,
    g1971_n
  );


  buf

  (
    g1972_n_spl_,
    g1972_n
  );


  buf

  (
    g1972_p_spl_,
    g1972_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    g1980_p_spl_,
    g1980_p
  );


  buf

  (
    g1981_p_spl_,
    g1981_p
  );


  buf

  (
    g1980_n_spl_,
    g1980_n
  );


  buf

  (
    g1981_n_spl_,
    g1981_n
  );


  buf

  (
    g1982_n_spl_,
    g1982_n
  );


  buf

  (
    g1982_n_spl_0,
    g1982_n_spl_
  );


  buf

  (
    g1982_p_spl_,
    g1982_p
  );


  buf

  (
    g1982_p_spl_0,
    g1982_p_spl_
  );


  buf

  (
    g1984_n_spl_,
    g1984_n
  );


  buf

  (
    g1984_p_spl_,
    g1984_p
  );


  buf

  (
    g1985_n_spl_,
    g1985_n
  );


  buf

  (
    g1985_p_spl_,
    g1985_p
  );


  buf

  (
    g1979_n_spl_,
    g1979_n
  );


  buf

  (
    g1987_p_spl_,
    g1987_p
  );


  buf

  (
    g1979_p_spl_,
    g1979_p
  );


  buf

  (
    g1987_n_spl_,
    g1987_n
  );


  buf

  (
    g1988_n_spl_,
    g1988_n
  );


  buf

  (
    g1988_p_spl_,
    g1988_p
  );


  buf

  (
    g1978_n_spl_,
    g1978_n
  );


  buf

  (
    g1990_p_spl_,
    g1990_p
  );


  buf

  (
    g1978_p_spl_,
    g1978_p
  );


  buf

  (
    g1990_n_spl_,
    g1990_n
  );


  buf

  (
    g1991_n_spl_,
    g1991_n
  );


  buf

  (
    g1991_p_spl_,
    g1991_p
  );


  buf

  (
    g1977_n_spl_,
    g1977_n
  );


  buf

  (
    g1993_p_spl_,
    g1993_p
  );


  buf

  (
    g1977_p_spl_,
    g1977_p
  );


  buf

  (
    g1993_n_spl_,
    g1993_n
  );


  buf

  (
    g1994_n_spl_,
    g1994_n
  );


  buf

  (
    g1994_p_spl_,
    g1994_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_01,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    g2002_p_spl_,
    g2002_p
  );


  buf

  (
    g2003_p_spl_,
    g2003_p
  );


  buf

  (
    g2002_n_spl_,
    g2002_n
  );


  buf

  (
    g2003_n_spl_,
    g2003_n
  );


  buf

  (
    g2004_n_spl_,
    g2004_n
  );


  buf

  (
    g2004_n_spl_0,
    g2004_n_spl_
  );


  buf

  (
    g2004_p_spl_,
    g2004_p
  );


  buf

  (
    g2004_p_spl_0,
    g2004_p_spl_
  );


  buf

  (
    g2006_n_spl_,
    g2006_n
  );


  buf

  (
    g2006_p_spl_,
    g2006_p
  );


  buf

  (
    g2007_n_spl_,
    g2007_n
  );


  buf

  (
    g2007_p_spl_,
    g2007_p
  );


  buf

  (
    g2001_n_spl_,
    g2001_n
  );


  buf

  (
    g2009_p_spl_,
    g2009_p
  );


  buf

  (
    g2001_p_spl_,
    g2001_p
  );


  buf

  (
    g2009_n_spl_,
    g2009_n
  );


  buf

  (
    g2010_n_spl_,
    g2010_n
  );


  buf

  (
    g2010_p_spl_,
    g2010_p
  );


  buf

  (
    g2000_n_spl_,
    g2000_n
  );


  buf

  (
    g2012_p_spl_,
    g2012_p
  );


  buf

  (
    g2000_p_spl_,
    g2000_p
  );


  buf

  (
    g2012_n_spl_,
    g2012_n
  );


  buf

  (
    g2013_n_spl_,
    g2013_n
  );


  buf

  (
    g2013_p_spl_,
    g2013_p
  );


  buf

  (
    g1999_n_spl_,
    g1999_n
  );


  buf

  (
    g2015_p_spl_,
    g2015_p
  );


  buf

  (
    g1999_p_spl_,
    g1999_p
  );


  buf

  (
    g2015_n_spl_,
    g2015_n
  );


  buf

  (
    g2016_n_spl_,
    g2016_n
  );


  buf

  (
    g2016_p_spl_,
    g2016_p
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_01,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    g2024_p_spl_,
    g2024_p
  );


  buf

  (
    g2025_p_spl_,
    g2025_p
  );


  buf

  (
    g2024_n_spl_,
    g2024_n
  );


  buf

  (
    g2025_n_spl_,
    g2025_n
  );


  buf

  (
    g2026_n_spl_,
    g2026_n
  );


  buf

  (
    g2026_n_spl_0,
    g2026_n_spl_
  );


  buf

  (
    g2026_p_spl_,
    g2026_p
  );


  buf

  (
    g2026_p_spl_0,
    g2026_p_spl_
  );


  buf

  (
    g2028_n_spl_,
    g2028_n
  );


  buf

  (
    g2028_p_spl_,
    g2028_p
  );


  buf

  (
    g2029_n_spl_,
    g2029_n
  );


  buf

  (
    g2029_p_spl_,
    g2029_p
  );


  buf

  (
    g2023_n_spl_,
    g2023_n
  );


  buf

  (
    g2031_p_spl_,
    g2031_p
  );


  buf

  (
    g2023_p_spl_,
    g2023_p
  );


  buf

  (
    g2031_n_spl_,
    g2031_n
  );


  buf

  (
    g2032_n_spl_,
    g2032_n
  );


  buf

  (
    g2032_p_spl_,
    g2032_p
  );


  buf

  (
    g2022_n_spl_,
    g2022_n
  );


  buf

  (
    g2034_p_spl_,
    g2034_p
  );


  buf

  (
    g2022_p_spl_,
    g2022_p
  );


  buf

  (
    g2034_n_spl_,
    g2034_n
  );


  buf

  (
    g2035_n_spl_,
    g2035_n
  );


  buf

  (
    g2035_p_spl_,
    g2035_p
  );


  buf

  (
    g2021_n_spl_,
    g2021_n
  );


  buf

  (
    g2037_p_spl_,
    g2037_p
  );


  buf

  (
    g2021_p_spl_,
    g2021_p
  );


  buf

  (
    g2037_n_spl_,
    g2037_n
  );


  buf

  (
    g2038_n_spl_,
    g2038_n
  );


  buf

  (
    g2038_p_spl_,
    g2038_p
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_01,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    g2046_p_spl_,
    g2046_p
  );


  buf

  (
    g2047_p_spl_,
    g2047_p
  );


  buf

  (
    g2046_n_spl_,
    g2046_n
  );


  buf

  (
    g2047_n_spl_,
    g2047_n
  );


  buf

  (
    g2048_n_spl_,
    g2048_n
  );


  buf

  (
    g2048_n_spl_0,
    g2048_n_spl_
  );


  buf

  (
    g2048_p_spl_,
    g2048_p
  );


  buf

  (
    g2048_p_spl_0,
    g2048_p_spl_
  );


  buf

  (
    g2050_n_spl_,
    g2050_n
  );


  buf

  (
    g2050_p_spl_,
    g2050_p
  );


  buf

  (
    g2051_n_spl_,
    g2051_n
  );


  buf

  (
    g2051_p_spl_,
    g2051_p
  );


  buf

  (
    g2045_n_spl_,
    g2045_n
  );


  buf

  (
    g2053_p_spl_,
    g2053_p
  );


  buf

  (
    g2045_p_spl_,
    g2045_p
  );


  buf

  (
    g2053_n_spl_,
    g2053_n
  );


  buf

  (
    g2054_n_spl_,
    g2054_n
  );


  buf

  (
    g2054_p_spl_,
    g2054_p
  );


  buf

  (
    g2044_n_spl_,
    g2044_n
  );


  buf

  (
    g2056_p_spl_,
    g2056_p
  );


  buf

  (
    g2044_p_spl_,
    g2044_p
  );


  buf

  (
    g2056_n_spl_,
    g2056_n
  );


  buf

  (
    g2057_n_spl_,
    g2057_n
  );


  buf

  (
    g2057_p_spl_,
    g2057_p
  );


  buf

  (
    g2043_n_spl_,
    g2043_n
  );


  buf

  (
    g2059_p_spl_,
    g2059_p
  );


  buf

  (
    g2043_p_spl_,
    g2043_p
  );


  buf

  (
    g2059_n_spl_,
    g2059_n
  );


  buf

  (
    g2060_n_spl_,
    g2060_n
  );


  buf

  (
    g2060_p_spl_,
    g2060_p
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    g2068_p_spl_,
    g2068_p
  );


  buf

  (
    g2069_p_spl_,
    g2069_p
  );


  buf

  (
    g2068_n_spl_,
    g2068_n
  );


  buf

  (
    g2069_n_spl_,
    g2069_n
  );


  buf

  (
    g2070_n_spl_,
    g2070_n
  );


  buf

  (
    g2070_n_spl_0,
    g2070_n_spl_
  );


  buf

  (
    g2070_p_spl_,
    g2070_p
  );


  buf

  (
    g2070_p_spl_0,
    g2070_p_spl_
  );


  buf

  (
    g2072_n_spl_,
    g2072_n
  );


  buf

  (
    g2072_p_spl_,
    g2072_p
  );


  buf

  (
    g2073_n_spl_,
    g2073_n
  );


  buf

  (
    g2073_p_spl_,
    g2073_p
  );


  buf

  (
    g2067_n_spl_,
    g2067_n
  );


  buf

  (
    g2075_p_spl_,
    g2075_p
  );


  buf

  (
    g2067_p_spl_,
    g2067_p
  );


  buf

  (
    g2075_n_spl_,
    g2075_n
  );


  buf

  (
    g2076_n_spl_,
    g2076_n
  );


  buf

  (
    g2076_p_spl_,
    g2076_p
  );


  buf

  (
    g2066_n_spl_,
    g2066_n
  );


  buf

  (
    g2078_p_spl_,
    g2078_p
  );


  buf

  (
    g2066_p_spl_,
    g2066_p
  );


  buf

  (
    g2078_n_spl_,
    g2078_n
  );


  buf

  (
    g2079_n_spl_,
    g2079_n
  );


  buf

  (
    g2079_p_spl_,
    g2079_p
  );


  buf

  (
    g2065_n_spl_,
    g2065_n
  );


  buf

  (
    g2081_p_spl_,
    g2081_p
  );


  buf

  (
    g2065_p_spl_,
    g2065_p
  );


  buf

  (
    g2081_n_spl_,
    g2081_n
  );


  buf

  (
    g2082_n_spl_,
    g2082_n
  );


  buf

  (
    g2082_p_spl_,
    g2082_p
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_01,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    g2090_p_spl_,
    g2090_p
  );


  buf

  (
    g2091_p_spl_,
    g2091_p
  );


  buf

  (
    g2090_n_spl_,
    g2090_n
  );


  buf

  (
    g2091_n_spl_,
    g2091_n
  );


  buf

  (
    g2092_n_spl_,
    g2092_n
  );


  buf

  (
    g2092_n_spl_0,
    g2092_n_spl_
  );


  buf

  (
    g2092_p_spl_,
    g2092_p
  );


  buf

  (
    g2092_p_spl_0,
    g2092_p_spl_
  );


  buf

  (
    g2094_n_spl_,
    g2094_n
  );


  buf

  (
    g2094_p_spl_,
    g2094_p
  );


  buf

  (
    g2095_n_spl_,
    g2095_n
  );


  buf

  (
    g2095_p_spl_,
    g2095_p
  );


  buf

  (
    g2089_n_spl_,
    g2089_n
  );


  buf

  (
    g2097_p_spl_,
    g2097_p
  );


  buf

  (
    g2089_p_spl_,
    g2089_p
  );


  buf

  (
    g2097_n_spl_,
    g2097_n
  );


  buf

  (
    g2098_n_spl_,
    g2098_n
  );


  buf

  (
    g2098_p_spl_,
    g2098_p
  );


  buf

  (
    g2088_n_spl_,
    g2088_n
  );


  buf

  (
    g2100_p_spl_,
    g2100_p
  );


  buf

  (
    g2088_p_spl_,
    g2088_p
  );


  buf

  (
    g2100_n_spl_,
    g2100_n
  );


  buf

  (
    g2101_n_spl_,
    g2101_n
  );


  buf

  (
    g2101_p_spl_,
    g2101_p
  );


  buf

  (
    g2087_n_spl_,
    g2087_n
  );


  buf

  (
    g2103_p_spl_,
    g2103_p
  );


  buf

  (
    g2087_p_spl_,
    g2087_p
  );


  buf

  (
    g2103_n_spl_,
    g2103_n
  );


  buf

  (
    g2104_n_spl_,
    g2104_n
  );


  buf

  (
    g2104_p_spl_,
    g2104_p
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_01,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    g2112_p_spl_,
    g2112_p
  );


  buf

  (
    g2113_p_spl_,
    g2113_p
  );


  buf

  (
    g2112_n_spl_,
    g2112_n
  );


  buf

  (
    g2113_n_spl_,
    g2113_n
  );


  buf

  (
    g2114_n_spl_,
    g2114_n
  );


  buf

  (
    g2114_n_spl_0,
    g2114_n_spl_
  );


  buf

  (
    g2114_p_spl_,
    g2114_p
  );


  buf

  (
    g2114_p_spl_0,
    g2114_p_spl_
  );


  buf

  (
    g2116_n_spl_,
    g2116_n
  );


  buf

  (
    g2116_p_spl_,
    g2116_p
  );


  buf

  (
    g2117_n_spl_,
    g2117_n
  );


  buf

  (
    g2117_p_spl_,
    g2117_p
  );


  buf

  (
    g2111_n_spl_,
    g2111_n
  );


  buf

  (
    g2119_p_spl_,
    g2119_p
  );


  buf

  (
    g2111_p_spl_,
    g2111_p
  );


  buf

  (
    g2119_n_spl_,
    g2119_n
  );


  buf

  (
    g2120_n_spl_,
    g2120_n
  );


  buf

  (
    g2120_p_spl_,
    g2120_p
  );


  buf

  (
    g2110_n_spl_,
    g2110_n
  );


  buf

  (
    g2122_p_spl_,
    g2122_p
  );


  buf

  (
    g2110_p_spl_,
    g2110_p
  );


  buf

  (
    g2122_n_spl_,
    g2122_n
  );


  buf

  (
    g2123_n_spl_,
    g2123_n
  );


  buf

  (
    g2123_p_spl_,
    g2123_p
  );


  buf

  (
    g2109_n_spl_,
    g2109_n
  );


  buf

  (
    g2125_p_spl_,
    g2125_p
  );


  buf

  (
    g2109_p_spl_,
    g2109_p
  );


  buf

  (
    g2125_n_spl_,
    g2125_n
  );


  buf

  (
    g2126_n_spl_,
    g2126_n
  );


  buf

  (
    g2126_p_spl_,
    g2126_p
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    g2134_p_spl_,
    g2134_p
  );


  buf

  (
    g2135_p_spl_,
    g2135_p
  );


  buf

  (
    g2134_n_spl_,
    g2134_n
  );


  buf

  (
    g2135_n_spl_,
    g2135_n
  );


  buf

  (
    g2136_n_spl_,
    g2136_n
  );


  buf

  (
    g2136_n_spl_0,
    g2136_n_spl_
  );


  buf

  (
    g2136_p_spl_,
    g2136_p
  );


  buf

  (
    g2136_p_spl_0,
    g2136_p_spl_
  );


  buf

  (
    g2138_n_spl_,
    g2138_n
  );


  buf

  (
    g2138_p_spl_,
    g2138_p
  );


  buf

  (
    g2139_n_spl_,
    g2139_n
  );


  buf

  (
    g2139_p_spl_,
    g2139_p
  );


  buf

  (
    g2133_n_spl_,
    g2133_n
  );


  buf

  (
    g2141_p_spl_,
    g2141_p
  );


  buf

  (
    g2133_p_spl_,
    g2133_p
  );


  buf

  (
    g2141_n_spl_,
    g2141_n
  );


  buf

  (
    g2142_n_spl_,
    g2142_n
  );


  buf

  (
    g2142_p_spl_,
    g2142_p
  );


  buf

  (
    g2132_n_spl_,
    g2132_n
  );


  buf

  (
    g2144_p_spl_,
    g2144_p
  );


  buf

  (
    g2132_p_spl_,
    g2132_p
  );


  buf

  (
    g2144_n_spl_,
    g2144_n
  );


  buf

  (
    g2145_n_spl_,
    g2145_n
  );


  buf

  (
    g2145_p_spl_,
    g2145_p
  );


  buf

  (
    g2131_n_spl_,
    g2131_n
  );


  buf

  (
    g2147_p_spl_,
    g2147_p
  );


  buf

  (
    g2131_p_spl_,
    g2131_p
  );


  buf

  (
    g2147_n_spl_,
    g2147_n
  );


  buf

  (
    g2148_n_spl_,
    g2148_n
  );


  buf

  (
    g2148_p_spl_,
    g2148_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    g2156_p_spl_,
    g2156_p
  );


  buf

  (
    g2157_p_spl_,
    g2157_p
  );


  buf

  (
    g2156_n_spl_,
    g2156_n
  );


  buf

  (
    g2157_n_spl_,
    g2157_n
  );


  buf

  (
    g2158_n_spl_,
    g2158_n
  );


  buf

  (
    g2158_p_spl_,
    g2158_p
  );


  buf

  (
    g2160_n_spl_,
    g2160_n
  );


  buf

  (
    g2160_p_spl_,
    g2160_p
  );


  buf

  (
    g2161_n_spl_,
    g2161_n
  );


  buf

  (
    g2161_p_spl_,
    g2161_p
  );


  buf

  (
    g2155_n_spl_,
    g2155_n
  );


  buf

  (
    g2163_p_spl_,
    g2163_p
  );


  buf

  (
    g2155_p_spl_,
    g2155_p
  );


  buf

  (
    g2163_n_spl_,
    g2163_n
  );


  buf

  (
    g2164_n_spl_,
    g2164_n
  );


  buf

  (
    g2164_p_spl_,
    g2164_p
  );


  buf

  (
    g2154_n_spl_,
    g2154_n
  );


  buf

  (
    g2166_p_spl_,
    g2166_p
  );


  buf

  (
    g2154_p_spl_,
    g2154_p
  );


  buf

  (
    g2166_n_spl_,
    g2166_n
  );


  buf

  (
    g2167_n_spl_,
    g2167_n
  );


  buf

  (
    g2167_p_spl_,
    g2167_p
  );


  buf

  (
    g2153_n_spl_,
    g2153_n
  );


  buf

  (
    g2169_p_spl_,
    g2169_p
  );


  buf

  (
    g2153_p_spl_,
    g2153_p
  );


  buf

  (
    g2169_n_spl_,
    g2169_n
  );


  buf

  (
    g2170_n_spl_,
    g2170_n
  );


  buf

  (
    g2170_p_spl_,
    g2170_p
  );


  buf

  (
    g2177_p_spl_,
    g2177_p
  );


  buf

  (
    g2177_n_spl_,
    g2177_n
  );


  buf

  (
    g2178_p_spl_,
    g2178_p
  );


  buf

  (
    g2179_n_spl_,
    g2179_n
  );


  buf

  (
    g2178_n_spl_,
    g2178_n
  );


  buf

  (
    g2179_p_spl_,
    g2179_p
  );


  buf

  (
    g2180_n_spl_,
    g2180_n
  );


  buf

  (
    g2180_p_spl_,
    g2180_p
  );


  buf

  (
    g2176_n_spl_,
    g2176_n
  );


  buf

  (
    g2182_p_spl_,
    g2182_p
  );


  buf

  (
    g2176_p_spl_,
    g2176_p
  );


  buf

  (
    g2182_n_spl_,
    g2182_n
  );


  buf

  (
    g2183_n_spl_,
    g2183_n
  );


  buf

  (
    g2183_p_spl_,
    g2183_p
  );


  buf

  (
    g2175_n_spl_,
    g2175_n
  );


  buf

  (
    g2185_p_spl_,
    g2185_p
  );


  buf

  (
    g2175_p_spl_,
    g2175_p
  );


  buf

  (
    g2185_n_spl_,
    g2185_n
  );


  buf

  (
    g2186_n_spl_,
    g2186_n
  );


  buf

  (
    g2186_p_spl_,
    g2186_p
  );


  buf

  (
    g2192_n_spl_,
    g2192_n
  );


  buf

  (
    g2193_n_spl_,
    g2193_n
  );


  buf

  (
    g2192_p_spl_,
    g2192_p
  );


  buf

  (
    g2193_p_spl_,
    g2193_p
  );


  buf

  (
    g2194_n_spl_,
    g2194_n
  );


  buf

  (
    g2191_n_spl_,
    g2191_n
  );


  buf

  (
    g2196_p_spl_,
    g2196_p
  );


  buf

  (
    g2191_p_spl_,
    g2191_p
  );


  buf

  (
    g2196_n_spl_,
    g2196_n
  );


  buf

  (
    g2197_n_spl_,
    g2197_n
  );


  buf

  (
    g2201_n_spl_,
    g2201_n
  );


  buf

  (
    g2203_p_spl_,
    g2203_p
  );


  buf

  (
    g2201_p_spl_,
    g2201_p
  );


  buf

  (
    g2203_n_spl_,
    g2203_n
  );


  buf

  (
    g2204_n_spl_,
    g2204_n
  );


  buf

  (
    g2204_p_spl_,
    g2204_p
  );


  buf

  (
    g2205_n_spl_,
    g2205_n
  );


  buf

  (
    g2207_p_spl_,
    g2207_p
  );


  buf

  (
    g2208_n_spl_,
    g2208_n
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_000,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_001,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_01,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_010,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_011,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_10,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_100,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_101,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_11,
    G21_p_spl_1
  );


  buf

  (
    g1631_p_spl_,
    g1631_p
  );


  buf

  (
    g2228_n_spl_,
    g2228_n
  );


  buf

  (
    g2230_p_spl_,
    g2230_p
  );


  buf

  (
    g1975_n_spl_,
    g1975_n
  );


  buf

  (
    g1997_n_spl_,
    g1997_n
  );


  buf

  (
    g2019_n_spl_,
    g2019_n
  );


  buf

  (
    g2041_n_spl_,
    g2041_n
  );


  buf

  (
    g2063_n_spl_,
    g2063_n
  );


  buf

  (
    g2085_n_spl_,
    g2085_n
  );


  buf

  (
    g2107_n_spl_,
    g2107_n
  );


  buf

  (
    g2129_n_spl_,
    g2129_n
  );


  buf

  (
    g2151_n_spl_,
    g2151_n
  );


  buf

  (
    g2173_n_spl_,
    g2173_n
  );


  buf

  (
    g2189_n_spl_,
    g2189_n
  );


  buf

  (
    g2200_n_spl_,
    g2200_n
  );


  buf

  (
    g2212_n_spl_,
    g2212_n
  );


endmodule
