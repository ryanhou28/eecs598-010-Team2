// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:58 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160,
    G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172,
    G173, G174, G175, G176, G177, G178,
    G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315;
  reg n2610_lo, n2613_lo, n2616_lo, n2619_lo, n2622_lo, n2625_lo, n2628_lo,
    n2631_lo, n2634_lo, n2637_lo, n2640_lo, n2643_lo, n2646_lo, n2649_lo,
    n2652_lo, n2655_lo, n2658_lo, n2661_lo, n2664_lo, n2667_lo, n2670_lo,
    n2673_lo, n2676_lo, n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo,
    n2694_lo, n2697_lo, n2700_lo, n2703_lo, n2706_lo, n2709_lo, n2712_lo,
    n2715_lo, n2718_lo, n2721_lo, n2724_lo, n2727_lo, n2730_lo, n2733_lo,
    n2736_lo, n2739_lo, n2742_lo, n2745_lo, n2748_lo, n2751_lo, n2754_lo,
    n2757_lo, n2760_lo, n2763_lo, n2766_lo, n2769_lo, n2772_lo, n2775_lo,
    n2778_lo, n2781_lo, n2784_lo, n2787_lo, n2790_lo, n2793_lo, n2796_lo,
    n2799_lo, n2802_lo, n2805_lo, n2808_lo, n2811_lo, n2814_lo, n2817_lo,
    n2820_lo, n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2835_lo, n2838_lo,
    n2841_lo, n2844_lo, n2847_lo, n2850_lo, n2853_lo, n2856_lo, n2859_lo,
    n2862_lo, n2865_lo, n2868_lo, n2871_lo, n2874_lo, n2877_lo, n2880_lo,
    n2883_lo, n2886_lo, n2889_lo, n2892_lo, n2895_lo, n2898_lo, n2901_lo,
    n2904_lo, n2907_lo, n2910_lo, n2913_lo, n2916_lo, n2919_lo, n2922_lo,
    n2925_lo, n2928_lo, n2931_lo, n2934_lo, n2937_lo, n2940_lo, n2943_lo,
    n2946_lo, n2949_lo, n2952_lo, n2955_lo, n2958_lo, n2961_lo, n2964_lo,
    n2967_lo, n2970_lo, n2973_lo, n2976_lo, n2979_lo, n2982_lo, n2985_lo,
    n2988_lo, n2991_lo, n2994_lo, n2997_lo, n3000_lo, n3003_lo, n3006_lo,
    n3009_lo, n3012_lo, n3015_lo, n3018_lo, n3021_lo, n3024_lo, n3027_lo,
    n3030_lo, n3033_lo, n3036_lo, n3039_lo, n3042_lo, n3045_lo, n3048_lo,
    n3051_lo, n3054_lo, n3057_lo, n3060_lo, n3063_lo, n3066_lo, n3069_lo,
    n3072_lo, n3075_lo, n3078_lo, n3081_lo, n3084_lo, n3087_lo, n3090_lo,
    n3093_lo, n3096_lo, n3099_lo, n3102_lo, n3105_lo, n3108_lo, n3111_lo,
    n3114_lo, n3117_lo, n3120_lo, n3123_lo, n3126_lo, n3129_lo, n3132_lo,
    n3135_lo, n3138_lo, n3141_lo, n3144_lo, n3147_lo, n3150_lo, n3153_lo,
    n3156_lo, n3159_lo, n3162_lo, n3165_lo, n3168_lo, n3171_lo, n3174_lo,
    n3177_lo, n3180_lo, n3183_lo, n3186_lo, n3189_lo, n3192_lo, n3195_lo,
    n3198_lo, n3201_lo, n3204_lo, n3207_lo, n3210_lo, n3213_lo, n3216_lo,
    n3219_lo, n3222_lo, n3225_lo, n3228_lo, n3231_lo, n3234_lo, n3237_lo,
    n3240_lo, n3243_lo, n3246_lo, n3249_lo, n3252_lo, n3255_lo, n3258_lo,
    n3261_lo, n3264_lo, n3267_lo, n3270_lo, n3273_lo, n3276_lo, n3279_lo,
    n3282_lo, n3285_lo, n3288_lo, n3291_lo, n3294_lo, n3297_lo, n3300_lo,
    n3303_lo, n3306_lo, n3309_lo, n3312_lo, n3315_lo, n3318_lo, n3321_lo,
    n3324_lo, n3327_lo, n3330_lo, n3333_lo, n3336_lo, n3339_lo, n3342_lo,
    n3345_lo, n3348_lo, n3351_lo, n3354_lo, n3357_lo, n3360_lo, n3363_lo,
    n3366_lo, n3369_lo, n3372_lo, n3375_lo, n3378_lo, n3381_lo, n3384_lo,
    n3387_lo, n3390_lo, n3393_lo, n3396_lo, n3399_lo, n3402_lo, n3405_lo,
    n3408_lo, n3411_lo, n3414_lo, n3417_lo, n3420_lo, n3423_lo, n3426_lo,
    n3429_lo, n3432_lo, n3435_lo, n3438_lo, n3441_lo, n3444_lo, n3447_lo,
    n3450_lo, n3453_lo, n3456_lo, n3459_lo, n3462_lo, n3465_lo, n3468_lo,
    n3471_lo, n3474_lo, n3477_lo, n3480_lo, n3483_lo, n3486_lo, n3489_lo,
    n3492_lo, n3495_lo, n3498_lo, n3501_lo, n3504_lo, n3507_lo, n3510_lo,
    n3513_lo, n3516_lo, n3519_lo, n3522_lo, n3525_lo, n3528_lo, n3531_lo,
    n3534_lo, n3537_lo, n3540_lo, n3543_lo, n3546_lo, n3549_lo, n3552_lo,
    n3555_lo, n3558_lo, n3561_lo, n3564_lo, n3567_lo, n3570_lo, n3573_lo,
    n3576_lo, n3579_lo, n3582_lo, n3585_lo, n3588_lo, n3591_lo, n3594_lo,
    n3597_lo, n3600_lo, n3603_lo, n3606_lo, n3609_lo, n3612_lo, n3615_lo,
    n3618_lo, n3621_lo, n3624_lo, n3627_lo, n3630_lo, n3633_lo, n3636_lo,
    n3639_lo, n3642_lo, n3645_lo, n3648_lo, n3651_lo, n3654_lo, n3657_lo,
    n3666_lo, n3669_lo, n3678_lo, n3687_lo, n3690_lo, n3702_lo, n3711_lo,
    n3714_lo, n3726_lo, n3735_lo, n3738_lo, n3750_lo, n3753_lo, n3759_lo,
    n3762_lo, n3765_lo, n3774_lo, n3777_lo, n3786_lo, n3789_lo, n3792_lo,
    n3795_lo, n3798_lo, n3801_lo, n3810_lo, n3813_lo, n3822_lo, n3825_lo,
    n3834_lo, n3843_lo, n3846_lo, n3867_lo, n3891_lo, n3915_lo, n3930_lo,
    n3933_lo, n3936_lo, n3942_lo, n3945_lo, n3948_lo, n3954_lo, n3957_lo,
    n3963_lo, n3966_lo, n3969_lo, n3975_lo, n3978_lo, n3987_lo, n3990_lo,
    n4002_lo, n4011_lo, n4014_lo, n4026_lo, n4035_lo, n4038_lo, n4050_lo,
    n4053_lo, n4059_lo, n4062_lo, n4065_lo, n4098_lo, n4107_lo, n4119_lo,
    n4131_lo, n4143_lo, n4155_lo, n4167_lo, n4179_lo, n4182_lo, n4185_lo,
    n4188_lo, n4194_lo, n4197_lo, n4200_lo, n4206_lo, n4209_lo, n4212_lo,
    n4215_lo, n4227_lo, n4230_lo, n4233_lo, n4236_lo, n4239_lo, n4242_lo,
    n4251_lo, n4263_lo, n4275_lo, n4278_lo, n4287_lo, n4290_lo, n4293_lo,
    n4299_lo, n4302_lo, n4305_lo, n4311_lo, n4314_lo, n4323_lo, n4326_lo,
    n4335_lo, n4338_lo, n4347_lo, n4350_lo, n4359_lo, n4362_lo, n4365_lo,
    n4371_lo, n4374_lo, n4383_lo, n4395_lo, n4407_lo, n4410_lo, n4413_lo,
    n4416_lo, n4419_lo, n4422_lo, n4425_lo, n4428_lo, n4431_lo, n4434_lo,
    n4437_lo, n4440_lo, n4443_lo, n4446_lo, n4449_lo, n4452_lo, n4455_lo,
    n4458_lo, n4461_lo, n4464_lo, n4467_lo, n4470_lo, n4473_lo, n4476_lo,
    n4479_lo, n4482_lo, n4485_lo, n4488_lo, n4494_lo, n4497_lo, n4500_lo,
    n4503_lo, n4506_lo, n4509_lo, n4512_lo, n4515_lo, n4518_lo, n4521_lo,
    n4524_lo, n4527_lo, n4530_lo, n4533_lo, n4536_lo, n4539_lo, n4542_lo,
    n4545_lo, n4548_lo, n4554_lo, n4557_lo, n4560_lo, n4563_lo, n4566_lo,
    n4569_lo, n4572_lo, n4575_lo, n4578_lo, n4581_lo, n4584_lo, n4587_lo,
    n4590_lo, n4593_lo, n4596_lo, n4599_lo, n4602_lo, n4605_lo, n4608_lo,
    n4611_lo, n4614_lo, n4617_lo, n4620_lo, n4623_lo, n4626_lo, n4629_lo,
    n4632_lo, n4635_lo, n4638_lo, n4641_lo, n4644_lo, n4647_lo, n4650_lo,
    n4653_lo, n4656_lo, n4659_lo, n4662_lo, n4665_lo, n4668_lo, n4671_lo,
    n4674_lo, n4677_lo, n4680_lo, n4683_lo, n4686_lo, n4689_lo, n4692_lo,
    n4695_lo, n4698_lo, n4701_lo, n4704_lo, n4707_lo, n4710_lo, n4713_lo,
    n4716_lo, n4719_lo, n4722_lo, n4725_lo, n4728_lo, n4731_lo, n4734_lo,
    n4737_lo, n4740_lo, n4743_lo, n6382_o2, n6383_o2, n6419_o2, n6420_o2,
    n6435_o2, n6436_o2, n6448_o2, n6449_o2, n6613_o2, n6614_o2, n6641_o2,
    n6658_o2, n6757_o2, n6756_o2, n7116_o2, n7156_o2, n6549_o2, n6550_o2,
    n7357_o2, n7358_o2, n7359_o2, n7360_o2, n6621_o2, n6623_o2, n6625_o2,
    n6626_o2, n6627_o2, n6628_o2, n6629_o2, n6630_o2, n6669_o2, n7449_o2,
    n7450_o2, n7451_o2, n7452_o2, n6682_o2, n6683_o2, n6684_o2, n6685_o2,
    n7463_o2, n6686_o2, n6687_o2, n6688_o2, n6689_o2, n6772_o2, n6773_o2,
    n6774_o2, n6775_o2, G3467_o2, G2810_o2, n6833_o2, n6945_o2, n6947_o2,
    n6949_o2, n6951_o2, n6888_o2, n6889_o2, n6936_o2, n6954_o2, n6955_o2,
    n6956_o2, n6957_o2, n6958_o2, n6982_o2, n6984_o2, n6974_o2, n6975_o2,
    n6999_o2, n7015_o2, n7016_o2, n7017_o2, n7018_o2, n7005_o2, n7019_o2,
    n7022_o2, n7023_o2, n7132_o2, n7133_o2, n7135_o2, n7136_o2, n7175_o2,
    n7155_o2, G3060_o2, n7383_o2, G3802_o2, G3859_o2, n7355_o2, n7356_o2,
    G4054_o2, G4068_o2, n7384_o2, n7387_o2, n7388_o2, n7389_o2, n7386_o2,
    n7453_o2, n7431_o2, n7432_o2, n7433_o2, n7430_o2, n7485_o2, n7486_o2,
    G2508_o2, G2486_o2, n2326_inv, n2329_inv, n3756_lo_buf_o2,
    n4056_lo_buf_o2, G3474_o2, n2341_inv, n7396_o2, n7398_o2, n7400_o2,
    n7401_o2, n7402_o2, n7403_o2, n7404_o2, n7405_o2, G2711_o2, n2371_inv,
    n7490_o2, n7527_o2, n7528_o2, n7529_o2, n7530_o2, n7523_o2, n7524_o2,
    n7525_o2, n7526_o2, n4296_lo_buf_o2, n4368_lo_buf_o2, G2466_o2,
    G2404_o2, n7534_o2, n7535_o2, n7536_o2, n7533_o2, G1060_o2, G963_o2,
    G2448_o2, G2685_o2, G2679_o2, G2774_o2, G2780_o2, G2759_o2, G2737_o2,
    G2850_o2, G3393_o2, G3404_o2, G3559_o2, G2744_o2, n3708_lo_buf_o2,
    n3840_lo_buf_o2, n4008_lo_buf_o2, n4104_lo_buf_o2, G1821_o2, G1734_o2,
    G3517_o2, G3533_o2, G3629_o2, G3645_o2, n2497_inv, G2731_o2, G2844_o2,
    n3732_lo_buf_o2, n4032_lo_buf_o2, G3552_o2, G2271_o2, n4248_lo_buf_o2,
    n4332_lo_buf_o2, n4344_lo_buf_o2, n4380_lo_buf_o2, G2398_o2, G2480_o2,
    G2418_o2, G1455_o2, G1449_o2, G1452_o2, G1425_o2, G1428_o2, G1419_o2,
    G1422_o2, n4308_lo_buf_o2, G2675_o2, G3035_o2, G3026_o2, G3029_o2,
    G3032_o2, G2999_o2, G3002_o2, G2770_o2, G3008_o2, G2073_o2, G2752_o2,
    G3005_o2, G5108_o2, G5135_o2, G5111_o2, G5138_o2, G3415_o2, G3386_o2,
    G3570_o2, G2430_o2, G3495_o2, G3621_o2, n4284_lo_buf_o2,
    n4356_lo_buf_o2, G2472_o2, G2410_o2, n3960_lo_buf_o2, n3972_lo_buf_o2,
    n2647_inv, n2650_inv, n3684_lo_buf_o2, n4080_lo_buf_o2,
    n4092_lo_buf_o2, n2662_inv, n2665_inv, G1147_o2, G2705_o2, G2693_o2,
    G2696_o2, G2700_o2, G2915_o2, G2966_o2, G2540_o2, G2788_o2, G2792_o2,
    G2797_o2, G2804_o2, G1038_o2, G1044_o2, G1090_o2, G1096_o2, G1029_o2,
    G3942_o2, G3954_o2, G4011_o2, G4017_o2, G1141_o2, G1081_o2, G2146_o2,
    G2145_o2, G2144_o2, G2143_o2, G2142_o2, G2141_o2, G2140_o2, G2139_o2,
    G3769_o2, G3773_o2, G3768_o2, G4101_o2, G3161_o2, G4143_o2, G3828_o2,
    G3831_o2, G3334_o2, G3335_o2, G3180_o2, G3340_o2, G3339_o2, G3341_o2,
    G3234_o2, G3829_o2, G3338_o2, G3336_o2, G3770_o2, G3918_o2, G3774_o2,
    G3921_o2, G3832_o2, G3993_o2, G2076_o2, G2071_o2, G2072_o2, G2069_o2,
    G2070_o2, G2067_o2, G2068_o2, G4095_o2, G3272_o2, G3269_o2, G3270_o2,
    G3271_o2, G3265_o2, G3266_o2, G4137_o2, G3268_o2, G2361_o2, G3228_o2,
    G3267_o2, G2336_o2, G3459_o2, G3428_o2, G3438_o2, G3449_o2, G3421_o2,
    G3576_o2, G3303_o2, G3583_o2, G3594_o2, G3674_o2, G3685_o2, G4504_o2,
    G4180_o2, G5123_o2, G5142_o2, G5126_o2, G5144_o2, G3912_o2, G4417_o2,
    G4420_o2, G3969_o2, G4023_o2, G2720_o2, G2837_o2, n2965_inv, n2968_inv,
    n2971_inv, n2974_inv, G1876_o2, G4996_o2, G4984_o2, G4920_o2, G4923_o2,
    G4930_o2, G4933_o2, n4320_lo_buf_o2, G2424_o2, G3317_o2, G3503_o2,
    G3485_o2, G3611_o2, n3864_lo_buf_o2, n3888_lo_buf_o2, n4116_lo_buf_o2,
    n4128_lo_buf_o2, n4140_lo_buf_o2, n4152_lo_buf_o2, G1815_o2, G1728_o2,
    G1035_o2, G1041_o2, G1087_o2, G1093_o2, G1132_o2, G1108_o2, G1138_o2,
    G1114_o2, G1807_o2, G2108_o2, G1126_o2, G1899_o2, G2134_o2, G1852_o2,
    G2116_o2, G2543_o2, G2727_o2, G2715_o2, G2832_o2, G1873_o2, G3291_o2,
    G5025_o2, G5036_o2, G3132_o2, G5038_o2, G5039_o2, n3118_inv, n3121_inv,
    n3124_inv, n3127_inv, n3984_lo_buf_o2, G1802_o2, G1804_o2, G1849_o2,
    G1851_o2, G2492_o2, G1799_o2, G4231_o2, G4234_o2, G4245_o2, G4247_o2,
    G1894_o2, G1846_o2, G4238_o2, G4249_o2, G2293_o2, G5022_o2, G5006_o2,
    G4944_o2, G4946_o2, G4954_o2, G4956_o2, G3546_o2, G3658_o2, G1344_o2,
    G2921_o2, n3912_lo_buf_o2, G1835_o2, G3810_o2, G3866_o2, G3811_o2,
    G2269_o2, G3812_o2, G3867_o2, G3868_o2, G3809_o2, G3716_o2, G4529_o2,
    G4670_o2, G4493_o2, G4580_o2, G3822_o2, G3877_o2, G4131_o2, G4170_o2,
    G4051_o2, G4065_o2, G4697_o2, G4706_o2, G2460_o2, G2454_o2, G2392_o2,
    G2386_o2, n4260_lo_buf_o2, n4272_lo_buf_o2, n4392_lo_buf_o2,
    n4404_lo_buf_o2, G1512_o2, G3135_o2, G2379_o2, n4164_lo_buf_o2,
    n4176_lo_buf_o2, n4224_lo_buf_o2, G2975_o2, G2978_o2, G2933_o2,
    G2936_o2, G1356_o2, G1359_o2, G1398_o2, G1401_o2;
  wire new_n2328_, new_n2330_, new_n2332_, new_n2334_, new_n2336_,
    new_n2338_, new_n2340_, new_n2342_, new_n2344_, new_n2346_, new_n2348_,
    new_n2350_, new_n2352_, new_n2354_, new_n2356_, new_n2358_, new_n2360_,
    new_n2362_, new_n2364_, new_n2366_, new_n2368_, new_n2370_, new_n2372_,
    new_n2374_, new_n2376_, new_n2378_, new_n2380_, new_n2382_, new_n2384_,
    new_n2386_, new_n2388_, new_n2390_, new_n2392_, new_n2394_, new_n2396_,
    new_n2398_, new_n2400_, new_n2402_, new_n2404_, new_n2406_, new_n2408_,
    new_n2410_, new_n2412_, new_n2414_, new_n2416_, new_n2418_, new_n2420_,
    new_n2422_, new_n2424_, new_n2426_, new_n2428_, new_n2430_, new_n2432_,
    new_n2434_, new_n2436_, new_n2438_, new_n2440_, new_n2442_, new_n2444_,
    new_n2446_, new_n2448_, new_n2450_, new_n2452_, new_n2454_, new_n2456_,
    new_n2458_, new_n2460_, new_n2462_, new_n2464_, new_n2466_, new_n2468_,
    new_n2470_, new_n2472_, new_n2474_, new_n2476_, new_n2478_, new_n2480_,
    new_n2482_, new_n2484_, new_n2486_, new_n2488_, new_n2490_, new_n2492_,
    new_n2494_, new_n2496_, new_n2498_, new_n2500_, new_n2502_, new_n2504_,
    new_n2506_, new_n2508_, new_n2510_, new_n2512_, new_n2514_, new_n2516_,
    new_n2518_, new_n2520_, new_n2522_, new_n2524_, new_n2526_, new_n2528_,
    new_n2530_, new_n2532_, new_n2534_, new_n2536_, new_n2538_, new_n2540_,
    new_n2542_, new_n2544_, new_n2546_, new_n2548_, new_n2550_, new_n2552_,
    new_n2554_, new_n2556_, new_n2558_, new_n2560_, new_n2562_, new_n2564_,
    new_n2566_, new_n2568_, new_n2570_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2578_, new_n2580_, new_n2582_, new_n2584_,
    new_n2586_, new_n2588_, new_n2590_, new_n2592_, new_n2594_, new_n2596_,
    new_n2598_, new_n2600_, new_n2602_, new_n2604_, new_n2606_, new_n2608_,
    new_n2610_, new_n2612_, new_n2614_, new_n2616_, new_n2618_, new_n2620_,
    new_n2622_, new_n2624_, new_n2626_, new_n2628_, new_n2630_, new_n2632_,
    new_n2634_, new_n2636_, new_n2638_, new_n2640_, new_n2642_, new_n2644_,
    new_n2646_, new_n2648_, new_n2650_, new_n2652_, new_n2654_, new_n2656_,
    new_n2658_, new_n2660_, new_n2662_, new_n2664_, new_n2666_, new_n2668_,
    new_n2670_, new_n2672_, new_n2674_, new_n2676_, new_n2678_, new_n2680_,
    new_n2682_, new_n2684_, new_n2686_, new_n2688_, new_n2690_, new_n2691_,
    new_n2692_, new_n2694_, new_n2696_, new_n2698_, new_n2699_, new_n2700_,
    new_n2702_, new_n2704_, new_n2706_, new_n2708_, new_n2710_, new_n2712_,
    new_n2714_, new_n2716_, new_n2718_, new_n2720_, new_n2722_, new_n2724_,
    new_n2726_, new_n2728_, new_n2730_, new_n2732_, new_n2734_, new_n2736_,
    new_n2739_, new_n2740_, new_n2742_, new_n2744_, new_n2747_, new_n2748_,
    new_n2750_, new_n2752_, new_n2755_, new_n2756_, new_n2758_, new_n2760_,
    new_n2763_, new_n2764_, new_n2766_, new_n2768_, new_n2770_, new_n2771_,
    new_n2772_, new_n2774_, new_n2776_, new_n2778_, new_n2779_, new_n2780_,
    new_n2782_, new_n2784_, new_n2787_, new_n2788_, new_n2790_, new_n2792_,
    new_n2794_, new_n2796_, new_n2798_, new_n2800_, new_n2802_, new_n2804_,
    new_n2806_, new_n2808_, new_n2810_, new_n2812_, new_n2814_, new_n2816_,
    new_n2818_, new_n2820_, new_n2822_, new_n2824_, new_n2826_, new_n2828_,
    new_n2830_, new_n2832_, new_n2834_, new_n2836_, new_n2838_, new_n2840_,
    new_n2842_, new_n2844_, new_n2846_, new_n2848_, new_n2850_, new_n2851_,
    new_n2852_, new_n2854_, new_n2856_, new_n2858_, new_n2860_, new_n2862_,
    new_n2864_, new_n2866_, new_n2868_, new_n2870_, new_n2872_, new_n2874_,
    new_n2876_, new_n2878_, new_n2880_, new_n2882_, new_n2884_, new_n2886_,
    new_n2888_, new_n2890_, new_n2892_, new_n2894_, new_n2896_, new_n2898_,
    new_n2900_, new_n2902_, new_n2904_, new_n2907_, new_n2908_, new_n2910_,
    new_n2912_, new_n2915_, new_n2916_, new_n2918_, new_n2920_, new_n2923_,
    new_n2924_, new_n2926_, new_n2928_, new_n2931_, new_n2932_, new_n2934_,
    new_n2936_, new_n2939_, new_n2940_, new_n2942_, new_n2944_, new_n2947_,
    new_n2948_, new_n2950_, new_n2952_, new_n2955_, new_n2956_, new_n2958_,
    new_n2960_, new_n2963_, new_n2964_, new_n2966_, new_n2968_, new_n2970_,
    new_n2972_, new_n2974_, new_n2976_, new_n2978_, new_n2980_, new_n2982_,
    new_n2984_, new_n2986_, new_n2988_, new_n2990_, new_n2992_, new_n2994_,
    new_n2996_, new_n2998_, new_n3000_, new_n3002_, new_n3004_, new_n3006_,
    new_n3008_, new_n3010_, new_n3012_, new_n3014_, new_n3016_, new_n3018_,
    new_n3020_, new_n3022_, new_n3024_, new_n3026_, new_n3028_, new_n3030_,
    new_n3032_, new_n3034_, new_n3036_, new_n3038_, new_n3040_, new_n3042_,
    new_n3044_, new_n3046_, new_n3048_, new_n3050_, new_n3052_, new_n3054_,
    new_n3056_, new_n3058_, new_n3060_, new_n3062_, new_n3064_, new_n3066_,
    new_n3068_, new_n3070_, new_n3072_, new_n3075_, new_n3076_, new_n3078_,
    new_n3080_, new_n3082_, new_n3084_, new_n3086_, new_n3088_, new_n3091_,
    new_n3092_, new_n3094_, new_n3096_, new_n3098_, new_n3100_, new_n3102_,
    new_n3104_, new_n3106_, new_n3108_, new_n3110_, new_n3112_, new_n3114_,
    new_n3116_, new_n3118_, new_n3120_, new_n3122_, new_n3124_, new_n3126_,
    new_n3128_, new_n3130_, new_n3132_, new_n3134_, new_n3136_, new_n3138_,
    new_n3140_, new_n3142_, new_n3144_, new_n3146_, new_n3148_, new_n3150_,
    new_n3152_, new_n3154_, new_n3156_, new_n3158_, new_n3160_, new_n3162_,
    new_n3164_, new_n3166_, new_n3168_, new_n3170_, new_n3171_, new_n3172_,
    new_n3174_, new_n3176_, new_n3179_, new_n3180_, new_n3182_, new_n3184_,
    new_n3186_, new_n3188_, new_n3190_, new_n3192_, new_n3194_, new_n3196_,
    new_n3198_, new_n3200_, new_n3203_, new_n3204_, new_n3206_, new_n3208_,
    new_n3210_, new_n3211_, new_n3212_, new_n3214_, new_n3216_, new_n3218_,
    new_n3220_, new_n3222_, new_n3224_, new_n3226_, new_n3228_, new_n3230_,
    new_n3232_, new_n3234_, new_n3236_, new_n3238_, new_n3240_, new_n3242_,
    new_n3244_, new_n3246_, new_n3248_, new_n3250_, new_n3252_, new_n3254_,
    new_n3256_, new_n3258_, new_n3260_, new_n3262_, new_n3264_, new_n3266_,
    new_n3268_, new_n3270_, new_n3272_, new_n3274_, new_n3276_, new_n3278_,
    new_n3280_, new_n3282_, new_n3284_, new_n3286_, new_n3288_, new_n3290_,
    new_n3292_, new_n3294_, new_n3296_, new_n3298_, new_n3300_, new_n3302_,
    new_n3304_, new_n3306_, new_n3308_, new_n3310_, new_n3312_, new_n3314_,
    new_n3316_, new_n3318_, new_n3320_, new_n3322_, new_n3324_, new_n3326_,
    new_n3328_, new_n3330_, new_n3332_, new_n3334_, new_n3336_, new_n3338_,
    new_n3340_, new_n3342_, new_n3344_, new_n3346_, new_n3348_, new_n3350_,
    new_n3352_, new_n3354_, new_n3356_, new_n3358_, new_n3360_, new_n3362_,
    new_n3364_, new_n3366_, new_n3368_, new_n3370_, new_n3372_, new_n3374_,
    new_n3376_, new_n3378_, new_n3380_, new_n3382_, new_n3384_, new_n3386_,
    new_n3388_, new_n3390_, new_n3391_, new_n3392_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3414_, new_n3415_,
    new_n3416_, new_n3418_, new_n3420_, new_n3422_, new_n3424_, new_n3427_,
    new_n3428_, new_n3430_, new_n3431_, new_n3432_, new_n3434_, new_n3435_,
    new_n3436_, new_n3438_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3454_, new_n3456_, new_n3457_,
    new_n3458_, new_n3460_, new_n3462_, new_n3463_, new_n3464_, new_n3466_,
    new_n3468_, new_n3469_, new_n3470_, new_n3472_, new_n3474_, new_n3475_,
    new_n3476_, new_n3478_, new_n3479_, new_n3480_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3507_, new_n3508_, new_n3509_, new_n3511_,
    new_n3512_, new_n3513_, new_n3515_, new_n3516_, new_n3517_, new_n3519_,
    new_n3520_, new_n3522_, new_n3524_, new_n3525_, new_n3526_, new_n3528_,
    new_n3530_, new_n3532_, new_n3534_, new_n3536_, new_n3538_, new_n3540_,
    new_n3541_, new_n3542_, new_n3544_, new_n3546_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3606_, new_n3608_, new_n3611_, new_n3612_,
    new_n3614_, new_n3616_, new_n3618_, new_n3619_, new_n3620_, new_n3622_,
    new_n3624_, new_n3626_, new_n3627_, new_n3628_, new_n3630_, new_n3632_,
    new_n3635_, new_n3636_, new_n3638_, new_n3640_, new_n3643_, new_n3644_,
    new_n3646_, new_n3648_, new_n3650_, new_n3651_, new_n3652_, new_n3654_,
    new_n3656_, new_n3657_, new_n3658_, new_n3660_, new_n3662_, new_n3664_,
    new_n3665_, new_n3666_, new_n3668_, new_n3670_, new_n3672_, new_n3673_,
    new_n3674_, new_n3676_, new_n3678_, new_n3680_, new_n3681_, new_n3682_,
    new_n3684_, new_n3686_, new_n3688_, new_n3689_, new_n3690_, new_n3692_,
    new_n3694_, new_n3695_, new_n3696_, new_n3698_, new_n3700_, new_n3702_,
    new_n3703_, new_n3704_, new_n3706_, new_n3708_, new_n3710_, new_n3712_,
    new_n3714_, new_n3716_, new_n3719_, new_n3720_, new_n3722_, new_n3724_,
    new_n3727_, new_n3728_, new_n3730_, new_n3732_, new_n3735_, new_n3736_,
    new_n3738_, new_n3740_, new_n3742_, new_n3744_, new_n3746_, new_n3748_,
    new_n3750_, new_n3752_, new_n3754_, new_n3756_, new_n3758_, new_n3759_,
    new_n3760_, new_n3762_, new_n3764_, new_n3766_, new_n3767_, new_n3768_,
    new_n3770_, new_n3772_, new_n3774_, new_n3775_, new_n3776_, new_n3778_,
    new_n3780_, new_n3782_, new_n3783_, new_n3784_, new_n3786_, new_n3788_,
    new_n3790_, new_n3791_, new_n3792_, new_n3794_, new_n3796_, new_n3798_,
    new_n3799_, new_n3800_, new_n3802_, new_n3804_, new_n3806_, new_n3807_,
    new_n3808_, new_n3810_, new_n3812_, new_n3814_, new_n3815_, new_n3816_,
    new_n3818_, new_n3820_, new_n3823_, new_n3825_, new_n3827_, new_n3829_,
    new_n3831_, new_n3833_, new_n3835_, new_n3837_, new_n3839_, new_n3841_,
    new_n3842_, new_n3845_, new_n3846_, new_n3848_, new_n3849_, new_n3850_,
    new_n3851_, new_n3853_, new_n3854_, new_n3855_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3862_, new_n3864_, new_n3866_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_,
    new_n3876_, new_n3877_, new_n3878_, new_n3880_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3889_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3916_,
    new_n3917_, new_n3918_, new_n3919_, new_n3921_, new_n3922_, new_n3924_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_,
    new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_,
    new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_,
    new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_,
    new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3989_, new_n3990_, new_n3991_, new_n3993_, new_n3995_,
    new_n3996_, new_n3998_, new_n4001_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4010_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4020_,
    new_n4022_, new_n4023_, new_n4024_, new_n4026_, new_n4028_, new_n4030_,
    new_n4031_, new_n4032_, new_n4034_, new_n4036_, new_n4037_, new_n4038_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4046_,
    new_n4048_, new_n4050_, new_n4052_, new_n4054_, new_n4056_, new_n4058_,
    new_n4060_, new_n4062_, new_n4064_, new_n4066_, new_n4068_, new_n4070_,
    new_n4072_, new_n4074_, new_n4076_, new_n4078_, new_n4080_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_,
    new_n4089_, new_n4090_, new_n4092_, new_n4094_, new_n4096_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4114_, new_n4116_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4126_,
    new_n4128_, new_n4129_, new_n4130_, new_n4132_, new_n4134_, new_n4135_,
    new_n4136_, new_n4137_, new_n4138_, new_n4140_, new_n4141_, new_n4142_,
    new_n4144_, new_n4145_, new_n4146_, new_n4148_, new_n4150_, new_n4152_,
    new_n4154_, new_n4156_, new_n4157_, new_n4158_, new_n4160_, new_n4162_,
    new_n4164_, new_n4166_, new_n4168_, new_n4170_, new_n4172_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4217_, new_n4219_,
    new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_,
    new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_,
    new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_,
    new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_,
    new_n4246_, new_n4247_, new_n4248_, new_n4250_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4437_, new_n4438_, new_n4440_, new_n4442_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4486_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4494_,
    new_n4496_, new_n4498_, new_n4500_, new_n4502_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_,
    new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_,
    new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_,
    new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_,
    new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_,
    new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n8443_, new_n8444_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_,
    new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_,
    new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_,
    new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_,
    new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_,
    new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_,
    new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_,
    new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_,
    new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_,
    new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_,
    new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_,
    new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_,
    new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_,
    new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_,
    new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_,
    new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_,
    new_n8878_, new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_,
    new_n8884_, new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_,
    new_n8890_, new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_,
    new_n8896_, new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_,
    new_n8914_, new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_,
    new_n8920_, new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_,
    new_n8926_, new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_,
    new_n8932_, new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_,
    new_n8938_, new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_,
    new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_,
    new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_,
    new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_,
    new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_,
    new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    n2610_li, n2613_li, n2616_li, n2619_li, n2622_li, n2625_li, n2628_li,
    n2631_li, n2634_li, n2637_li, n2640_li, n2643_li, n2646_li, n2649_li,
    n2652_li, n2655_li, n2658_li, n2661_li, n2664_li, n2667_li, n2670_li,
    n2673_li, n2676_li, n2679_li, n2682_li, n2685_li, n2688_li, n2691_li,
    n2694_li, n2697_li, n2700_li, n2703_li, n2706_li, n2709_li, n2712_li,
    n2715_li, n2718_li, n2721_li, n2724_li, n2727_li, n2730_li, n2733_li,
    n2736_li, n2739_li, n2742_li, n2745_li, n2748_li, n2751_li, n2754_li,
    n2757_li, n2760_li, n2763_li, n2766_li, n2769_li, n2772_li, n2775_li,
    n2778_li, n2781_li, n2784_li, n2787_li, n2790_li, n2793_li, n2796_li,
    n2799_li, n2802_li, n2805_li, n2808_li, n2811_li, n2814_li, n2817_li,
    n2820_li, n2823_li, n2826_li, n2829_li, n2832_li, n2835_li, n2838_li,
    n2841_li, n2844_li, n2847_li, n2850_li, n2853_li, n2856_li, n2859_li,
    n2862_li, n2865_li, n2868_li, n2871_li, n2874_li, n2877_li, n2880_li,
    n2883_li, n2886_li, n2889_li, n2892_li, n2895_li, n2898_li, n2901_li,
    n2904_li, n2907_li, n2910_li, n2913_li, n2916_li, n2919_li, n2922_li,
    n2925_li, n2928_li, n2931_li, n2934_li, n2937_li, n2940_li, n2943_li,
    n2946_li, n2949_li, n2952_li, n2955_li, n2958_li, n2961_li, n2964_li,
    n2967_li, n2970_li, n2973_li, n2976_li, n2979_li, n2982_li, n2985_li,
    n2988_li, n2991_li, n2994_li, n2997_li, n3000_li, n3003_li, n3006_li,
    n3009_li, n3012_li, n3015_li, n3018_li, n3021_li, n3024_li, n3027_li,
    n3030_li, n3033_li, n3036_li, n3039_li, n3042_li, n3045_li, n3048_li,
    n3051_li, n3054_li, n3057_li, n3060_li, n3063_li, n3066_li, n3069_li,
    n3072_li, n3075_li, n3078_li, n3081_li, n3084_li, n3087_li, n3090_li,
    n3093_li, n3096_li, n3099_li, n3102_li, n3105_li, n3108_li, n3111_li,
    n3114_li, n3117_li, n3120_li, n3123_li, n3126_li, n3129_li, n3132_li,
    n3135_li, n3138_li, n3141_li, n3144_li, n3147_li, n3150_li, n3153_li,
    n3156_li, n3159_li, n3162_li, n3165_li, n3168_li, n3171_li, n3174_li,
    n3177_li, n3180_li, n3183_li, n3186_li, n3189_li, n3192_li, n3195_li,
    n3198_li, n3201_li, n3204_li, n3207_li, n3210_li, n3213_li, n3216_li,
    n3219_li, n3222_li, n3225_li, n3228_li, n3231_li, n3234_li, n3237_li,
    n3240_li, n3243_li, n3246_li, n3249_li, n3252_li, n3255_li, n3258_li,
    n3261_li, n3264_li, n3267_li, n3270_li, n3273_li, n3276_li, n3279_li,
    n3282_li, n3285_li, n3288_li, n3291_li, n3294_li, n3297_li, n3300_li,
    n3303_li, n3306_li, n3309_li, n3312_li, n3315_li, n3318_li, n3321_li,
    n3324_li, n3327_li, n3330_li, n3333_li, n3336_li, n3339_li, n3342_li,
    n3345_li, n3348_li, n3351_li, n3354_li, n3357_li, n3360_li, n3363_li,
    n3366_li, n3369_li, n3372_li, n3375_li, n3378_li, n3381_li, n3384_li,
    n3387_li, n3390_li, n3393_li, n3396_li, n3399_li, n3402_li, n3405_li,
    n3408_li, n3411_li, n3414_li, n3417_li, n3420_li, n3423_li, n3426_li,
    n3429_li, n3432_li, n3435_li, n3438_li, n3441_li, n3444_li, n3447_li,
    n3450_li, n3453_li, n3456_li, n3459_li, n3462_li, n3465_li, n3468_li,
    n3471_li, n3474_li, n3477_li, n3480_li, n3483_li, n3486_li, n3489_li,
    n3492_li, n3495_li, n3498_li, n3501_li, n3504_li, n3507_li, n3510_li,
    n3513_li, n3516_li, n3519_li, n3522_li, n3525_li, n3528_li, n3531_li,
    n3534_li, n3537_li, n3540_li, n3543_li, n3546_li, n3549_li, n3552_li,
    n3555_li, n3558_li, n3561_li, n3564_li, n3567_li, n3570_li, n3573_li,
    n3576_li, n3579_li, n3582_li, n3585_li, n3588_li, n3591_li, n3594_li,
    n3597_li, n3600_li, n3603_li, n3606_li, n3609_li, n3612_li, n3615_li,
    n3618_li, n3621_li, n3624_li, n3627_li, n3630_li, n3633_li, n3636_li,
    n3639_li, n3642_li, n3645_li, n3648_li, n3651_li, n3654_li, n3657_li,
    n3666_li, n3669_li, n3678_li, n3687_li, n3690_li, n3702_li, n3711_li,
    n3714_li, n3726_li, n3735_li, n3738_li, n3750_li, n3753_li, n3759_li,
    n3762_li, n3765_li, n3774_li, n3777_li, n3786_li, n3789_li, n3792_li,
    n3795_li, n3798_li, n3801_li, n3810_li, n3813_li, n3822_li, n3825_li,
    n3834_li, n3843_li, n3846_li, n3867_li, n3891_li, n3915_li, n3930_li,
    n3933_li, n3936_li, n3942_li, n3945_li, n3948_li, n3954_li, n3957_li,
    n3963_li, n3966_li, n3969_li, n3975_li, n3978_li, n3987_li, n3990_li,
    n4002_li, n4011_li, n4014_li, n4026_li, n4035_li, n4038_li, n4050_li,
    n4053_li, n4059_li, n4062_li, n4065_li, n4098_li, n4107_li, n4119_li,
    n4131_li, n4143_li, n4155_li, n4167_li, n4179_li, n4182_li, n4185_li,
    n4188_li, n4194_li, n4197_li, n4200_li, n4206_li, n4209_li, n4212_li,
    n4215_li, n4227_li, n4230_li, n4233_li, n4236_li, n4239_li, n4242_li,
    n4251_li, n4263_li, n4275_li, n4278_li, n4287_li, n4290_li, n4293_li,
    n4299_li, n4302_li, n4305_li, n4311_li, n4314_li, n4323_li, n4326_li,
    n4335_li, n4338_li, n4347_li, n4350_li, n4359_li, n4362_li, n4365_li,
    n4371_li, n4374_li, n4383_li, n4395_li, n4407_li, n4410_li, n4413_li,
    n4416_li, n4419_li, n4422_li, n4425_li, n4428_li, n4431_li, n4434_li,
    n4437_li, n4440_li, n4443_li, n4446_li, n4449_li, n4452_li, n4455_li,
    n4458_li, n4461_li, n4464_li, n4467_li, n4470_li, n4473_li, n4476_li,
    n4479_li, n4482_li, n4485_li, n4488_li, n4494_li, n4497_li, n4500_li,
    n4503_li, n4506_li, n4509_li, n4512_li, n4515_li, n4518_li, n4521_li,
    n4524_li, n4527_li, n4530_li, n4533_li, n4536_li, n4539_li, n4542_li,
    n4545_li, n4548_li, n4554_li, n4557_li, n4560_li, n4563_li, n4566_li,
    n4569_li, n4572_li, n4575_li, n4578_li, n4581_li, n4584_li, n4587_li,
    n4590_li, n4593_li, n4596_li, n4599_li, n4602_li, n4605_li, n4608_li,
    n4611_li, n4614_li, n4617_li, n4620_li, n4623_li, n4626_li, n4629_li,
    n4632_li, n4635_li, n4638_li, n4641_li, n4644_li, n4647_li, n4650_li,
    n4653_li, n4656_li, n4659_li, n4662_li, n4665_li, n4668_li, n4671_li,
    n4674_li, n4677_li, n4680_li, n4683_li, n4686_li, n4689_li, n4692_li,
    n4695_li, n4698_li, n4701_li, n4704_li, n4707_li, n4710_li, n4713_li,
    n4716_li, n4719_li, n4722_li, n4725_li, n4728_li, n4731_li, n4734_li,
    n4737_li, n4740_li, n4743_li, n6382_i2, n6383_i2, n6419_i2, n6420_i2,
    n6435_i2, n6436_i2, n6448_i2, n6449_i2, n6613_i2, n6614_i2, n6641_i2,
    n6658_i2, n6757_i2, n6756_i2, n7116_i2, n7156_i2, n6549_i2, n6550_i2,
    n7357_i2, n7358_i2, n7359_i2, n7360_i2, n6621_i2, n6623_i2, n6625_i2,
    n6626_i2, n6627_i2, n6628_i2, n6629_i2, n6630_i2, n6669_i2, n7449_i2,
    n7450_i2, n7451_i2, n7452_i2, n6682_i2, n6683_i2, n6684_i2, n6685_i2,
    n7463_i2, n6686_i2, n6687_i2, n6688_i2, n6689_i2, n6772_i2, n6773_i2,
    n6774_i2, n6775_i2, G3467_i2, G2810_i2, n6833_i2, n6945_i2, n6947_i2,
    n6949_i2, n6951_i2, n6888_i2, n6889_i2, n6936_i2, n6954_i2, n6955_i2,
    n6956_i2, n6957_i2, n6958_i2, n6982_i2, n6984_i2, n6974_i2, n6975_i2,
    n6999_i2, n7015_i2, n7016_i2, n7017_i2, n7018_i2, n7005_i2, n7019_i2,
    n7022_i2, n7023_i2, n7132_i2, n7133_i2, n7135_i2, n7136_i2, n7175_i2,
    n7155_i2, G3060_i2, n7383_i2, G3802_i2, G3859_i2, n7355_i2, n7356_i2,
    G4054_i2, G4068_i2, n7384_i2, n7387_i2, n7388_i2, n7389_i2, n7386_i2,
    n7453_i2, n7431_i2, n7432_i2, n7433_i2, n7430_i2, n7485_i2, n7486_i2,
    G2508_i2, G2486_i2, n7245_i2, n7246_i2, n3756_lo_buf_i2,
    n4056_lo_buf_i2, G3474_i2, G2817_i2, n7396_i2, n7398_i2, n7400_i2,
    n7401_i2, n7402_i2, n7403_i2, n7404_i2, n7405_i2, G2711_i2, G2828_i2,
    n7490_i2, n7527_i2, n7528_i2, n7529_i2, n7530_i2, n7523_i2, n7524_i2,
    n7525_i2, n7526_i2, n4296_lo_buf_i2, n4368_lo_buf_i2, G2466_i2,
    G2404_i2, n7534_i2, n7535_i2, n7536_i2, n7533_i2, G1060_i2, G963_i2,
    G2448_i2, G2685_i2, G2679_i2, G2774_i2, G2780_i2, G2759_i2, G2737_i2,
    G2850_i2, G3393_i2, G3404_i2, G3559_i2, G2744_i2, n3708_lo_buf_i2,
    n3840_lo_buf_i2, n4008_lo_buf_i2, n4104_lo_buf_i2, G1821_i2, G1734_i2,
    G3517_i2, G3533_i2, G3629_i2, G3645_i2, G2857_i2, G2731_i2, G2844_i2,
    n3732_lo_buf_i2, n4032_lo_buf_i2, G3552_i2, G2271_i2, n4248_lo_buf_i2,
    n4332_lo_buf_i2, n4344_lo_buf_i2, n4380_lo_buf_i2, G2398_i2, G2480_i2,
    G2418_i2, G1455_i2, G1449_i2, G1452_i2, G1425_i2, G1428_i2, G1419_i2,
    G1422_i2, n4308_lo_buf_i2, G2675_i2, G3035_i2, G3026_i2, G3029_i2,
    G3032_i2, G2999_i2, G3002_i2, G2770_i2, G3008_i2, G2073_i2, G2752_i2,
    G3005_i2, G5108_i2, G5135_i2, G5111_i2, G5138_i2, G3415_i2, G3386_i2,
    G3570_i2, G2430_i2, G3495_i2, G3621_i2, n4284_lo_buf_i2,
    n4356_lo_buf_i2, G2472_i2, G2410_i2, n3960_lo_buf_i2, n3972_lo_buf_i2,
    G2865_i2, G970_i2, n3684_lo_buf_i2, n4080_lo_buf_i2, n4092_lo_buf_i2,
    G1053_i2, G956_i2, G1147_i2, G2705_i2, G2693_i2, G2696_i2, G2700_i2,
    G2915_i2, G2966_i2, G2540_i2, G2788_i2, G2792_i2, G2797_i2, G2804_i2,
    G1038_i2, G1044_i2, G1090_i2, G1096_i2, G1029_i2, G3942_i2, G3954_i2,
    G4011_i2, G4017_i2, G1141_i2, G1081_i2, G2146_i2, G2145_i2, G2144_i2,
    G2143_i2, G2142_i2, G2141_i2, G2140_i2, G2139_i2, G3769_i2, G3773_i2,
    G3768_i2, G4101_i2, G3161_i2, G4143_i2, G3828_i2, G3831_i2, G3334_i2,
    G3335_i2, G3180_i2, G3340_i2, G3339_i2, G3341_i2, G3234_i2, G3829_i2,
    G3338_i2, G3336_i2, G3770_i2, G3918_i2, G3774_i2, G3921_i2, G3832_i2,
    G3993_i2, G2076_i2, G2071_i2, G2072_i2, G2069_i2, G2070_i2, G2067_i2,
    G2068_i2, G4095_i2, G3272_i2, G3269_i2, G3270_i2, G3271_i2, G3265_i2,
    G3266_i2, G4137_i2, G3268_i2, G2361_i2, G3228_i2, G3267_i2, G2336_i2,
    G3459_i2, G3428_i2, G3438_i2, G3449_i2, G3421_i2, G3576_i2, G3303_i2,
    G3583_i2, G3594_i2, G3674_i2, G3685_i2, G4504_i2, G4180_i2, G5123_i2,
    G5142_i2, G5126_i2, G5144_i2, G3912_i2, G4417_i2, G4420_i2, G3969_i2,
    G4023_i2, G2720_i2, G2837_i2, G836_i2, G848_i2, G813_i2, G825_i2,
    G1876_i2, G4996_i2, G4984_i2, G4920_i2, G4923_i2, G4930_i2, G4933_i2,
    n4320_lo_buf_i2, G2424_i2, G3317_i2, G3503_i2, G3485_i2, G3611_i2,
    n3864_lo_buf_i2, n3888_lo_buf_i2, n4116_lo_buf_i2, n4128_lo_buf_i2,
    n4140_lo_buf_i2, n4152_lo_buf_i2, G1815_i2, G1728_i2, G1035_i2,
    G1041_i2, G1087_i2, G1093_i2, G1132_i2, G1108_i2, G1138_i2, G1114_i2,
    G1807_i2, G2108_i2, G1126_i2, G1899_i2, G2134_i2, G1852_i2, G2116_i2,
    G2543_i2, G2727_i2, G2715_i2, G2832_i2, G1873_i2, G3291_i2, G5025_i2,
    G5036_i2, G3132_i2, G5038_i2, G5039_i2, G1150_i2, G1162_i2, G804_i2,
    G1172_i2, n3984_lo_buf_i2, G1802_i2, G1804_i2, G1849_i2, G1851_i2,
    G2492_i2, G1799_i2, G4231_i2, G4234_i2, G4245_i2, G4247_i2, G1894_i2,
    G1846_i2, G4238_i2, G4249_i2, G2293_i2, G5022_i2, G5006_i2, G4944_i2,
    G4946_i2, G4954_i2, G4956_i2, G3546_i2, G3658_i2, G1344_i2, G2921_i2,
    n3912_lo_buf_i2, G1835_i2, G3810_i2, G3866_i2, G3811_i2, G2269_i2,
    G3812_i2, G3867_i2, G3868_i2, G3809_i2, G3716_i2, G4529_i2, G4670_i2,
    G4493_i2, G4580_i2, G3822_i2, G3877_i2, G4131_i2, G4170_i2, G4051_i2,
    G4065_i2, G4697_i2, G4706_i2, G2460_i2, G2454_i2, G2392_i2, G2386_i2,
    n4260_lo_buf_i2, n4272_lo_buf_i2, n4392_lo_buf_i2, n4404_lo_buf_i2,
    G1512_i2, G3135_i2, G2379_i2, n4164_lo_buf_i2, n4176_lo_buf_i2,
    n4224_lo_buf_i2, G2975_i2, G2978_i2, G2933_i2, G2936_i2, G1356_i2,
    G1359_i2, G1398_i2, G1401_i2;
  assign new_n2328_ = G1;
  assign new_n2330_ = G2;
  assign new_n2332_ = G3;
  assign new_n2334_ = G4;
  assign new_n2336_ = G5;
  assign new_n2338_ = G6;
  assign new_n2340_ = G7;
  assign new_n2342_ = G8;
  assign new_n2344_ = G9;
  assign new_n2346_ = G10;
  assign new_n2348_ = G11;
  assign new_n2350_ = G12;
  assign new_n2352_ = G13;
  assign new_n2354_ = G14;
  assign new_n2356_ = G15;
  assign new_n2358_ = G16;
  assign new_n2360_ = G17;
  assign new_n2362_ = G18;
  assign new_n2364_ = G19;
  assign new_n2366_ = G20;
  assign new_n2368_ = G21;
  assign new_n2370_ = G22;
  assign new_n2372_ = G23;
  assign new_n2374_ = G24;
  assign new_n2376_ = G25;
  assign new_n2378_ = G26;
  assign new_n2380_ = G27;
  assign new_n2382_ = G28;
  assign new_n2384_ = G29;
  assign new_n2386_ = G30;
  assign new_n2388_ = G31;
  assign new_n2390_ = G32;
  assign new_n2392_ = G33;
  assign new_n2394_ = G34;
  assign new_n2396_ = G35;
  assign new_n2398_ = G36;
  assign new_n2400_ = G37;
  assign new_n2402_ = G38;
  assign new_n2404_ = G39;
  assign new_n2406_ = G40;
  assign new_n2408_ = G41;
  assign new_n2410_ = G42;
  assign new_n2412_ = G43;
  assign new_n2414_ = G44;
  assign new_n2416_ = G45;
  assign new_n2418_ = G46;
  assign new_n2420_ = G47;
  assign new_n2422_ = G48;
  assign new_n2424_ = G49;
  assign new_n2426_ = G50;
  assign new_n2428_ = G51;
  assign new_n2430_ = G52;
  assign new_n2432_ = G53;
  assign new_n2434_ = G54;
  assign new_n2436_ = G55;
  assign new_n2438_ = G56;
  assign new_n2440_ = G57;
  assign new_n2442_ = G58;
  assign new_n2444_ = G59;
  assign new_n2446_ = G60;
  assign new_n2448_ = G61;
  assign new_n2450_ = G62;
  assign new_n2452_ = G63;
  assign new_n2454_ = G64;
  assign new_n2456_ = G65;
  assign new_n2458_ = G66;
  assign new_n2460_ = G67;
  assign new_n2462_ = G68;
  assign new_n2464_ = G69;
  assign new_n2466_ = G70;
  assign new_n2468_ = G71;
  assign new_n2470_ = G72;
  assign new_n2472_ = G73;
  assign new_n2474_ = G74;
  assign new_n2476_ = G75;
  assign new_n2478_ = G76;
  assign new_n2480_ = G77;
  assign new_n2482_ = G78;
  assign new_n2484_ = G79;
  assign new_n2486_ = G80;
  assign new_n2488_ = G81;
  assign new_n2490_ = G82;
  assign new_n2492_ = G83;
  assign new_n2494_ = G84;
  assign new_n2496_ = G85;
  assign new_n2498_ = G86;
  assign new_n2500_ = G87;
  assign new_n2502_ = G88;
  assign new_n2504_ = G89;
  assign new_n2506_ = G90;
  assign new_n2508_ = G91;
  assign new_n2510_ = G92;
  assign new_n2512_ = G93;
  assign new_n2514_ = G94;
  assign new_n2516_ = G95;
  assign new_n2518_ = G96;
  assign new_n2520_ = G97;
  assign new_n2522_ = G98;
  assign new_n2524_ = G99;
  assign new_n2526_ = G100;
  assign new_n2528_ = G101;
  assign new_n2530_ = G102;
  assign new_n2532_ = G103;
  assign new_n2534_ = G104;
  assign new_n2536_ = G105;
  assign new_n2538_ = G106;
  assign new_n2540_ = G107;
  assign new_n2542_ = G108;
  assign new_n2544_ = G109;
  assign new_n2546_ = G110;
  assign new_n2548_ = G111;
  assign new_n2550_ = G112;
  assign new_n2552_ = G113;
  assign new_n2554_ = G114;
  assign new_n2556_ = G115;
  assign new_n2558_ = G116;
  assign new_n2560_ = G117;
  assign new_n2562_ = G118;
  assign new_n2564_ = G119;
  assign new_n2566_ = G120;
  assign new_n2568_ = G121;
  assign new_n2570_ = G122;
  assign new_n2572_ = G123;
  assign new_n2573_ = ~G123;
  assign new_n2574_ = G124;
  assign new_n2575_ = ~G124;
  assign new_n2576_ = G125;
  assign new_n2578_ = G126;
  assign new_n2580_ = G127;
  assign new_n2582_ = G128;
  assign new_n2584_ = G129;
  assign new_n2586_ = G130;
  assign new_n2588_ = G131;
  assign new_n2590_ = G132;
  assign new_n2592_ = G133;
  assign new_n2594_ = G134;
  assign new_n2596_ = G135;
  assign new_n2598_ = G136;
  assign new_n2600_ = G137;
  assign new_n2602_ = G138;
  assign new_n2604_ = G139;
  assign new_n2606_ = G140;
  assign new_n2608_ = G141;
  assign new_n2610_ = G142;
  assign new_n2612_ = G143;
  assign new_n2614_ = G144;
  assign new_n2616_ = G145;
  assign new_n2618_ = G146;
  assign new_n2620_ = G147;
  assign new_n2622_ = G148;
  assign new_n2624_ = G149;
  assign new_n2626_ = G150;
  assign new_n2628_ = G151;
  assign new_n2630_ = G152;
  assign new_n2632_ = G153;
  assign new_n2634_ = G154;
  assign new_n2636_ = G155;
  assign new_n2638_ = G156;
  assign new_n2640_ = G157;
  assign new_n2642_ = G158;
  assign new_n2644_ = G159;
  assign new_n2646_ = G160;
  assign new_n2648_ = G161;
  assign new_n2650_ = G162;
  assign new_n2652_ = G163;
  assign new_n2654_ = G164;
  assign new_n2656_ = G165;
  assign new_n2658_ = G166;
  assign new_n2660_ = G167;
  assign new_n2662_ = G168;
  assign new_n2664_ = G169;
  assign new_n2666_ = G170;
  assign new_n2668_ = G171;
  assign new_n2670_ = G172;
  assign new_n2672_ = G173;
  assign new_n2674_ = G174;
  assign new_n2676_ = G175;
  assign new_n2678_ = G176;
  assign new_n2680_ = G177;
  assign new_n2682_ = G178;
  assign new_n2684_ = n2610_lo;
  assign new_n2686_ = n2613_lo;
  assign new_n2688_ = n2616_lo;
  assign new_n2690_ = n2619_lo;
  assign new_n2691_ = ~n2619_lo;
  assign new_n2692_ = n2622_lo;
  assign new_n2694_ = n2625_lo;
  assign new_n2696_ = n2628_lo;
  assign new_n2698_ = n2631_lo;
  assign new_n2699_ = ~n2631_lo;
  assign new_n2700_ = n2634_lo;
  assign new_n2702_ = n2637_lo;
  assign new_n2704_ = n2640_lo;
  assign new_n2706_ = n2643_lo;
  assign new_n2708_ = n2646_lo;
  assign new_n2710_ = n2649_lo;
  assign new_n2712_ = n2652_lo;
  assign new_n2714_ = n2655_lo;
  assign new_n2716_ = n2658_lo;
  assign new_n2718_ = n2661_lo;
  assign new_n2720_ = n2664_lo;
  assign new_n2722_ = n2667_lo;
  assign new_n2724_ = n2670_lo;
  assign new_n2726_ = n2673_lo;
  assign new_n2728_ = n2676_lo;
  assign new_n2730_ = n2679_lo;
  assign new_n2732_ = n2682_lo;
  assign new_n2734_ = n2685_lo;
  assign new_n2736_ = n2688_lo;
  assign new_n2739_ = ~n2691_lo;
  assign new_n2740_ = n2694_lo;
  assign new_n2742_ = n2697_lo;
  assign new_n2744_ = n2700_lo;
  assign new_n2747_ = ~n2703_lo;
  assign new_n2748_ = n2706_lo;
  assign new_n2750_ = n2709_lo;
  assign new_n2752_ = n2712_lo;
  assign new_n2755_ = ~n2715_lo;
  assign new_n2756_ = n2718_lo;
  assign new_n2758_ = n2721_lo;
  assign new_n2760_ = n2724_lo;
  assign new_n2763_ = ~n2727_lo;
  assign new_n2764_ = n2730_lo;
  assign new_n2766_ = n2733_lo;
  assign new_n2768_ = n2736_lo;
  assign new_n2770_ = n2739_lo;
  assign new_n2771_ = ~n2739_lo;
  assign new_n2772_ = n2742_lo;
  assign new_n2774_ = n2745_lo;
  assign new_n2776_ = n2748_lo;
  assign new_n2778_ = n2751_lo;
  assign new_n2779_ = ~n2751_lo;
  assign new_n2780_ = n2754_lo;
  assign new_n2782_ = n2757_lo;
  assign new_n2784_ = n2760_lo;
  assign new_n2787_ = ~n2763_lo;
  assign new_n2788_ = n2766_lo;
  assign new_n2790_ = n2769_lo;
  assign new_n2792_ = n2772_lo;
  assign new_n2794_ = n2775_lo;
  assign new_n2796_ = n2778_lo;
  assign new_n2798_ = n2781_lo;
  assign new_n2800_ = n2784_lo;
  assign new_n2802_ = n2787_lo;
  assign new_n2804_ = n2790_lo;
  assign new_n2806_ = n2793_lo;
  assign new_n2808_ = n2796_lo;
  assign new_n2810_ = n2799_lo;
  assign new_n2812_ = n2802_lo;
  assign new_n2814_ = n2805_lo;
  assign new_n2816_ = n2808_lo;
  assign new_n2818_ = n2811_lo;
  assign new_n2820_ = n2814_lo;
  assign new_n2822_ = n2817_lo;
  assign new_n2824_ = n2820_lo;
  assign new_n2826_ = n2823_lo;
  assign new_n2828_ = n2826_lo;
  assign new_n2830_ = n2829_lo;
  assign new_n2832_ = n2832_lo;
  assign new_n2834_ = n2835_lo;
  assign new_n2836_ = n2838_lo;
  assign new_n2838_ = n2841_lo;
  assign new_n2840_ = n2844_lo;
  assign new_n2842_ = n2847_lo;
  assign new_n2844_ = n2850_lo;
  assign new_n2846_ = n2853_lo;
  assign new_n2848_ = n2856_lo;
  assign new_n2850_ = n2859_lo;
  assign new_n2851_ = ~n2859_lo;
  assign new_n2852_ = n2862_lo;
  assign new_n2854_ = n2865_lo;
  assign new_n2856_ = n2868_lo;
  assign new_n2858_ = n2871_lo;
  assign new_n2860_ = n2874_lo;
  assign new_n2862_ = n2877_lo;
  assign new_n2864_ = n2880_lo;
  assign new_n2866_ = n2883_lo;
  assign new_n2868_ = n2886_lo;
  assign new_n2870_ = n2889_lo;
  assign new_n2872_ = n2892_lo;
  assign new_n2874_ = n2895_lo;
  assign new_n2876_ = n2898_lo;
  assign new_n2878_ = n2901_lo;
  assign new_n2880_ = n2904_lo;
  assign new_n2882_ = n2907_lo;
  assign new_n2884_ = n2910_lo;
  assign new_n2886_ = n2913_lo;
  assign new_n2888_ = n2916_lo;
  assign new_n2890_ = n2919_lo;
  assign new_n2892_ = n2922_lo;
  assign new_n2894_ = n2925_lo;
  assign new_n2896_ = n2928_lo;
  assign new_n2898_ = n2931_lo;
  assign new_n2900_ = n2934_lo;
  assign new_n2902_ = n2937_lo;
  assign new_n2904_ = n2940_lo;
  assign new_n2907_ = ~n2943_lo;
  assign new_n2908_ = n2946_lo;
  assign new_n2910_ = n2949_lo;
  assign new_n2912_ = n2952_lo;
  assign new_n2915_ = ~n2955_lo;
  assign new_n2916_ = n2958_lo;
  assign new_n2918_ = n2961_lo;
  assign new_n2920_ = n2964_lo;
  assign new_n2923_ = ~n2967_lo;
  assign new_n2924_ = n2970_lo;
  assign new_n2926_ = n2973_lo;
  assign new_n2928_ = n2976_lo;
  assign new_n2931_ = ~n2979_lo;
  assign new_n2932_ = n2982_lo;
  assign new_n2934_ = n2985_lo;
  assign new_n2936_ = n2988_lo;
  assign new_n2939_ = ~n2991_lo;
  assign new_n2940_ = n2994_lo;
  assign new_n2942_ = n2997_lo;
  assign new_n2944_ = n3000_lo;
  assign new_n2947_ = ~n3003_lo;
  assign new_n2948_ = n3006_lo;
  assign new_n2950_ = n3009_lo;
  assign new_n2952_ = n3012_lo;
  assign new_n2955_ = ~n3015_lo;
  assign new_n2956_ = n3018_lo;
  assign new_n2958_ = n3021_lo;
  assign new_n2960_ = n3024_lo;
  assign new_n2963_ = ~n3027_lo;
  assign new_n2964_ = n3030_lo;
  assign new_n2966_ = n3033_lo;
  assign new_n2968_ = n3036_lo;
  assign new_n2970_ = n3039_lo;
  assign new_n2972_ = n3042_lo;
  assign new_n2974_ = n3045_lo;
  assign new_n2976_ = n3048_lo;
  assign new_n2978_ = n3051_lo;
  assign new_n2980_ = n3054_lo;
  assign new_n2982_ = n3057_lo;
  assign new_n2984_ = n3060_lo;
  assign new_n2986_ = n3063_lo;
  assign new_n2988_ = n3066_lo;
  assign new_n2990_ = n3069_lo;
  assign new_n2992_ = n3072_lo;
  assign new_n2994_ = n3075_lo;
  assign new_n2996_ = n3078_lo;
  assign new_n2998_ = n3081_lo;
  assign new_n3000_ = n3084_lo;
  assign new_n3002_ = n3087_lo;
  assign new_n3004_ = n3090_lo;
  assign new_n3006_ = n3093_lo;
  assign new_n3008_ = n3096_lo;
  assign new_n3010_ = n3099_lo;
  assign new_n3012_ = n3102_lo;
  assign new_n3014_ = n3105_lo;
  assign new_n3016_ = n3108_lo;
  assign new_n3018_ = n3111_lo;
  assign new_n3020_ = n3114_lo;
  assign new_n3022_ = n3117_lo;
  assign new_n3024_ = n3120_lo;
  assign new_n3026_ = n3123_lo;
  assign new_n3028_ = n3126_lo;
  assign new_n3030_ = n3129_lo;
  assign new_n3032_ = n3132_lo;
  assign new_n3034_ = n3135_lo;
  assign new_n3036_ = n3138_lo;
  assign new_n3038_ = n3141_lo;
  assign new_n3040_ = n3144_lo;
  assign new_n3042_ = n3147_lo;
  assign new_n3044_ = n3150_lo;
  assign new_n3046_ = n3153_lo;
  assign new_n3048_ = n3156_lo;
  assign new_n3050_ = n3159_lo;
  assign new_n3052_ = n3162_lo;
  assign new_n3054_ = n3165_lo;
  assign new_n3056_ = n3168_lo;
  assign new_n3058_ = n3171_lo;
  assign new_n3060_ = n3174_lo;
  assign new_n3062_ = n3177_lo;
  assign new_n3064_ = n3180_lo;
  assign new_n3066_ = n3183_lo;
  assign new_n3068_ = n3186_lo;
  assign new_n3070_ = n3189_lo;
  assign new_n3072_ = n3192_lo;
  assign new_n3075_ = ~n3195_lo;
  assign new_n3076_ = n3198_lo;
  assign new_n3078_ = n3201_lo;
  assign new_n3080_ = n3204_lo;
  assign new_n3082_ = n3207_lo;
  assign new_n3084_ = n3210_lo;
  assign new_n3086_ = n3213_lo;
  assign new_n3088_ = n3216_lo;
  assign new_n3091_ = ~n3219_lo;
  assign new_n3092_ = n3222_lo;
  assign new_n3094_ = n3225_lo;
  assign new_n3096_ = n3228_lo;
  assign new_n3098_ = n3231_lo;
  assign new_n3100_ = n3234_lo;
  assign new_n3102_ = n3237_lo;
  assign new_n3104_ = n3240_lo;
  assign new_n3106_ = n3243_lo;
  assign new_n3108_ = n3246_lo;
  assign new_n3110_ = n3249_lo;
  assign new_n3112_ = n3252_lo;
  assign new_n3114_ = n3255_lo;
  assign new_n3116_ = n3258_lo;
  assign new_n3118_ = n3261_lo;
  assign new_n3120_ = n3264_lo;
  assign new_n3122_ = n3267_lo;
  assign new_n3124_ = n3270_lo;
  assign new_n3126_ = n3273_lo;
  assign new_n3128_ = n3276_lo;
  assign new_n3130_ = n3279_lo;
  assign new_n3132_ = n3282_lo;
  assign new_n3134_ = n3285_lo;
  assign new_n3136_ = n3288_lo;
  assign new_n3138_ = n3291_lo;
  assign new_n3140_ = n3294_lo;
  assign new_n3142_ = n3297_lo;
  assign new_n3144_ = n3300_lo;
  assign new_n3146_ = n3303_lo;
  assign new_n3148_ = n3306_lo;
  assign new_n3150_ = n3309_lo;
  assign new_n3152_ = n3312_lo;
  assign new_n3154_ = n3315_lo;
  assign new_n3156_ = n3318_lo;
  assign new_n3158_ = n3321_lo;
  assign new_n3160_ = n3324_lo;
  assign new_n3162_ = n3327_lo;
  assign new_n3164_ = n3330_lo;
  assign new_n3166_ = n3333_lo;
  assign new_n3168_ = n3336_lo;
  assign new_n3170_ = n3339_lo;
  assign new_n3171_ = ~n3339_lo;
  assign new_n3172_ = n3342_lo;
  assign new_n3174_ = n3345_lo;
  assign new_n3176_ = n3348_lo;
  assign new_n3179_ = ~n3351_lo;
  assign new_n3180_ = n3354_lo;
  assign new_n3182_ = n3357_lo;
  assign new_n3184_ = n3360_lo;
  assign new_n3186_ = n3363_lo;
  assign new_n3188_ = n3366_lo;
  assign new_n3190_ = n3369_lo;
  assign new_n3192_ = n3372_lo;
  assign new_n3194_ = n3375_lo;
  assign new_n3196_ = n3378_lo;
  assign new_n3198_ = n3381_lo;
  assign new_n3200_ = n3384_lo;
  assign new_n3203_ = ~n3387_lo;
  assign new_n3204_ = n3390_lo;
  assign new_n3206_ = n3393_lo;
  assign new_n3208_ = n3396_lo;
  assign new_n3210_ = n3399_lo;
  assign new_n3211_ = ~n3399_lo;
  assign new_n3212_ = n3402_lo;
  assign new_n3214_ = n3405_lo;
  assign new_n3216_ = n3408_lo;
  assign new_n3218_ = n3411_lo;
  assign new_n3220_ = n3414_lo;
  assign new_n3222_ = n3417_lo;
  assign new_n3224_ = n3420_lo;
  assign new_n3226_ = n3423_lo;
  assign new_n3228_ = n3426_lo;
  assign new_n3230_ = n3429_lo;
  assign new_n3232_ = n3432_lo;
  assign new_n3234_ = n3435_lo;
  assign new_n3236_ = n3438_lo;
  assign new_n3238_ = n3441_lo;
  assign new_n3240_ = n3444_lo;
  assign new_n3242_ = n3447_lo;
  assign new_n3244_ = n3450_lo;
  assign new_n3246_ = n3453_lo;
  assign new_n3248_ = n3456_lo;
  assign new_n3250_ = n3459_lo;
  assign new_n3252_ = n3462_lo;
  assign new_n3254_ = n3465_lo;
  assign new_n3256_ = n3468_lo;
  assign new_n3258_ = n3471_lo;
  assign new_n3260_ = n3474_lo;
  assign new_n3262_ = n3477_lo;
  assign new_n3264_ = n3480_lo;
  assign new_n3266_ = n3483_lo;
  assign new_n3268_ = n3486_lo;
  assign new_n3270_ = n3489_lo;
  assign new_n3272_ = n3492_lo;
  assign new_n3274_ = n3495_lo;
  assign new_n3276_ = n3498_lo;
  assign new_n3278_ = n3501_lo;
  assign new_n3280_ = n3504_lo;
  assign new_n3282_ = n3507_lo;
  assign new_n3284_ = n3510_lo;
  assign new_n3286_ = n3513_lo;
  assign new_n3288_ = n3516_lo;
  assign new_n3290_ = n3519_lo;
  assign new_n3292_ = n3522_lo;
  assign new_n3294_ = n3525_lo;
  assign new_n3296_ = n3528_lo;
  assign new_n3298_ = n3531_lo;
  assign new_n3300_ = n3534_lo;
  assign new_n3302_ = n3537_lo;
  assign new_n3304_ = n3540_lo;
  assign new_n3306_ = n3543_lo;
  assign new_n3308_ = n3546_lo;
  assign new_n3310_ = n3549_lo;
  assign new_n3312_ = n3552_lo;
  assign new_n3314_ = n3555_lo;
  assign new_n3316_ = n3558_lo;
  assign new_n3318_ = n3561_lo;
  assign new_n3320_ = n3564_lo;
  assign new_n3322_ = n3567_lo;
  assign new_n3324_ = n3570_lo;
  assign new_n3326_ = n3573_lo;
  assign new_n3328_ = n3576_lo;
  assign new_n3330_ = n3579_lo;
  assign new_n3332_ = n3582_lo;
  assign new_n3334_ = n3585_lo;
  assign new_n3336_ = n3588_lo;
  assign new_n3338_ = n3591_lo;
  assign new_n3340_ = n3594_lo;
  assign new_n3342_ = n3597_lo;
  assign new_n3344_ = n3600_lo;
  assign new_n3346_ = n3603_lo;
  assign new_n3348_ = n3606_lo;
  assign new_n3350_ = n3609_lo;
  assign new_n3352_ = n3612_lo;
  assign new_n3354_ = n3615_lo;
  assign new_n3356_ = n3618_lo;
  assign new_n3358_ = n3621_lo;
  assign new_n3360_ = n3624_lo;
  assign new_n3362_ = n3627_lo;
  assign new_n3364_ = n3630_lo;
  assign new_n3366_ = n3633_lo;
  assign new_n3368_ = n3636_lo;
  assign new_n3370_ = n3639_lo;
  assign new_n3372_ = n3642_lo;
  assign new_n3374_ = n3645_lo;
  assign new_n3376_ = n3648_lo;
  assign new_n3378_ = n3651_lo;
  assign new_n3380_ = n3654_lo;
  assign new_n3382_ = n3657_lo;
  assign new_n3384_ = n3666_lo;
  assign new_n3386_ = n3669_lo;
  assign new_n3388_ = n3678_lo;
  assign new_n3390_ = n3687_lo;
  assign new_n3391_ = ~n3687_lo;
  assign new_n3392_ = n3690_lo;
  assign new_n3394_ = n3702_lo;
  assign new_n3395_ = ~n3702_lo;
  assign new_n3396_ = n3711_lo;
  assign new_n3397_ = ~n3711_lo;
  assign new_n3398_ = n3714_lo;
  assign new_n3399_ = ~n3714_lo;
  assign new_n3400_ = n3726_lo;
  assign new_n3401_ = ~n3726_lo;
  assign new_n3402_ = n3735_lo;
  assign new_n3403_ = ~n3735_lo;
  assign new_n3404_ = n3738_lo;
  assign new_n3405_ = ~n3738_lo;
  assign new_n3406_ = n3750_lo;
  assign new_n3408_ = n3753_lo;
  assign new_n3409_ = ~n3753_lo;
  assign new_n3410_ = n3759_lo;
  assign new_n3411_ = ~n3759_lo;
  assign new_n3412_ = n3762_lo;
  assign new_n3414_ = n3765_lo;
  assign new_n3415_ = ~n3765_lo;
  assign new_n3416_ = n3774_lo;
  assign new_n3418_ = n3777_lo;
  assign new_n3420_ = n3786_lo;
  assign new_n3422_ = n3789_lo;
  assign new_n3424_ = n3792_lo;
  assign new_n3427_ = ~n3795_lo;
  assign new_n3428_ = n3798_lo;
  assign new_n3430_ = n3801_lo;
  assign new_n3431_ = ~n3801_lo;
  assign new_n3432_ = n3810_lo;
  assign new_n3434_ = n3813_lo;
  assign new_n3435_ = ~n3813_lo;
  assign new_n3436_ = n3822_lo;
  assign new_n3438_ = n3825_lo;
  assign new_n3440_ = n3834_lo;
  assign new_n3441_ = ~n3834_lo;
  assign new_n3442_ = n3843_lo;
  assign new_n3443_ = ~n3843_lo;
  assign new_n3444_ = n3846_lo;
  assign new_n3445_ = ~n3846_lo;
  assign new_n3446_ = n3867_lo;
  assign new_n3447_ = ~n3867_lo;
  assign new_n3448_ = n3891_lo;
  assign new_n3449_ = ~n3891_lo;
  assign new_n3450_ = n3915_lo;
  assign new_n3451_ = ~n3915_lo;
  assign new_n3452_ = n3930_lo;
  assign new_n3454_ = n3933_lo;
  assign new_n3456_ = n3936_lo;
  assign new_n3457_ = ~n3936_lo;
  assign new_n3458_ = n3942_lo;
  assign new_n3460_ = n3945_lo;
  assign new_n3462_ = n3948_lo;
  assign new_n3463_ = ~n3948_lo;
  assign new_n3464_ = n3954_lo;
  assign new_n3466_ = n3957_lo;
  assign new_n3468_ = n3963_lo;
  assign new_n3469_ = ~n3963_lo;
  assign new_n3470_ = n3966_lo;
  assign new_n3472_ = n3969_lo;
  assign new_n3474_ = n3975_lo;
  assign new_n3475_ = ~n3975_lo;
  assign new_n3476_ = n3978_lo;
  assign new_n3478_ = n3987_lo;
  assign new_n3479_ = ~n3987_lo;
  assign new_n3480_ = n3990_lo;
  assign new_n3482_ = n4002_lo;
  assign new_n3483_ = ~n4002_lo;
  assign new_n3484_ = n4011_lo;
  assign new_n3485_ = ~n4011_lo;
  assign new_n3486_ = n4014_lo;
  assign new_n3487_ = ~n4014_lo;
  assign new_n3488_ = n4026_lo;
  assign new_n3489_ = ~n4026_lo;
  assign new_n3490_ = n4035_lo;
  assign new_n3491_ = ~n4035_lo;
  assign new_n3492_ = n4038_lo;
  assign new_n3493_ = ~n4038_lo;
  assign new_n3494_ = n4050_lo;
  assign new_n3496_ = n4053_lo;
  assign new_n3497_ = ~n4053_lo;
  assign new_n3498_ = n4059_lo;
  assign new_n3499_ = ~n4059_lo;
  assign new_n3500_ = n4062_lo;
  assign new_n3502_ = n4065_lo;
  assign new_n3503_ = ~n4065_lo;
  assign new_n3504_ = n4098_lo;
  assign new_n3505_ = ~n4098_lo;
  assign new_n3507_ = ~n4107_lo;
  assign new_n3508_ = n4119_lo;
  assign new_n3509_ = ~n4119_lo;
  assign new_n3511_ = ~n4131_lo;
  assign new_n3512_ = n4143_lo;
  assign new_n3513_ = ~n4143_lo;
  assign new_n3515_ = ~n4155_lo;
  assign new_n3516_ = n4167_lo;
  assign new_n3517_ = ~n4167_lo;
  assign new_n3519_ = ~n4179_lo;
  assign new_n3520_ = n4182_lo;
  assign new_n3522_ = n4185_lo;
  assign new_n3524_ = n4188_lo;
  assign new_n3525_ = ~n4188_lo;
  assign new_n3526_ = n4194_lo;
  assign new_n3528_ = n4197_lo;
  assign new_n3530_ = n4200_lo;
  assign new_n3532_ = n4206_lo;
  assign new_n3534_ = n4209_lo;
  assign new_n3536_ = n4212_lo;
  assign new_n3538_ = n4215_lo;
  assign new_n3540_ = n4227_lo;
  assign new_n3541_ = ~n4227_lo;
  assign new_n3542_ = n4230_lo;
  assign new_n3544_ = n4233_lo;
  assign new_n3546_ = n4236_lo;
  assign new_n3549_ = ~n4239_lo;
  assign new_n3550_ = n4242_lo;
  assign new_n3551_ = ~n4242_lo;
  assign new_n3552_ = n4251_lo;
  assign new_n3553_ = ~n4251_lo;
  assign new_n3554_ = n4263_lo;
  assign new_n3555_ = ~n4263_lo;
  assign new_n3556_ = n4275_lo;
  assign new_n3557_ = ~n4275_lo;
  assign new_n3558_ = n4278_lo;
  assign new_n3559_ = ~n4278_lo;
  assign new_n3560_ = n4287_lo;
  assign new_n3561_ = ~n4287_lo;
  assign new_n3562_ = n4290_lo;
  assign new_n3564_ = n4293_lo;
  assign new_n3565_ = ~n4293_lo;
  assign new_n3566_ = n4299_lo;
  assign new_n3567_ = ~n4299_lo;
  assign new_n3568_ = n4302_lo;
  assign new_n3570_ = n4305_lo;
  assign new_n3571_ = ~n4305_lo;
  assign new_n3572_ = n4311_lo;
  assign new_n3573_ = ~n4311_lo;
  assign new_n3574_ = n4314_lo;
  assign new_n3576_ = n4323_lo;
  assign new_n3577_ = ~n4323_lo;
  assign new_n3578_ = n4326_lo;
  assign new_n3579_ = ~n4326_lo;
  assign new_n3580_ = n4335_lo;
  assign new_n3581_ = ~n4335_lo;
  assign new_n3582_ = n4338_lo;
  assign new_n3583_ = ~n4338_lo;
  assign new_n3584_ = n4347_lo;
  assign new_n3585_ = ~n4347_lo;
  assign new_n3586_ = n4350_lo;
  assign new_n3587_ = ~n4350_lo;
  assign new_n3588_ = n4359_lo;
  assign new_n3589_ = ~n4359_lo;
  assign new_n3590_ = n4362_lo;
  assign new_n3592_ = n4365_lo;
  assign new_n3593_ = ~n4365_lo;
  assign new_n3594_ = n4371_lo;
  assign new_n3595_ = ~n4371_lo;
  assign new_n3596_ = n4374_lo;
  assign new_n3597_ = ~n4374_lo;
  assign new_n3598_ = n4383_lo;
  assign new_n3599_ = ~n4383_lo;
  assign new_n3600_ = n4395_lo;
  assign new_n3601_ = ~n4395_lo;
  assign new_n3602_ = n4407_lo;
  assign new_n3603_ = ~n4407_lo;
  assign new_n3604_ = n4410_lo;
  assign new_n3606_ = n4413_lo;
  assign new_n3608_ = n4416_lo;
  assign new_n3611_ = ~n4419_lo;
  assign new_n3612_ = n4422_lo;
  assign new_n3614_ = n4425_lo;
  assign new_n3616_ = n4428_lo;
  assign new_n3618_ = n4431_lo;
  assign new_n3619_ = ~n4431_lo;
  assign new_n3620_ = n4434_lo;
  assign new_n3622_ = n4437_lo;
  assign new_n3624_ = n4440_lo;
  assign new_n3626_ = n4443_lo;
  assign new_n3627_ = ~n4443_lo;
  assign new_n3628_ = n4446_lo;
  assign new_n3630_ = n4449_lo;
  assign new_n3632_ = n4452_lo;
  assign new_n3635_ = ~n4455_lo;
  assign new_n3636_ = n4458_lo;
  assign new_n3638_ = n4461_lo;
  assign new_n3640_ = n4464_lo;
  assign new_n3643_ = ~n4467_lo;
  assign new_n3644_ = n4470_lo;
  assign new_n3646_ = n4473_lo;
  assign new_n3648_ = n4476_lo;
  assign new_n3650_ = n4479_lo;
  assign new_n3651_ = ~n4479_lo;
  assign new_n3652_ = n4482_lo;
  assign new_n3654_ = n4485_lo;
  assign new_n3656_ = n4488_lo;
  assign new_n3657_ = ~n4488_lo;
  assign new_n3658_ = n4494_lo;
  assign new_n3660_ = n4497_lo;
  assign new_n3662_ = n4500_lo;
  assign new_n3664_ = n4503_lo;
  assign new_n3665_ = ~n4503_lo;
  assign new_n3666_ = n4506_lo;
  assign new_n3668_ = n4509_lo;
  assign new_n3670_ = n4512_lo;
  assign new_n3672_ = n4515_lo;
  assign new_n3673_ = ~n4515_lo;
  assign new_n3674_ = n4518_lo;
  assign new_n3676_ = n4521_lo;
  assign new_n3678_ = n4524_lo;
  assign new_n3680_ = n4527_lo;
  assign new_n3681_ = ~n4527_lo;
  assign new_n3682_ = n4530_lo;
  assign new_n3684_ = n4533_lo;
  assign new_n3686_ = n4536_lo;
  assign new_n3688_ = n4539_lo;
  assign new_n3689_ = ~n4539_lo;
  assign new_n3690_ = n4542_lo;
  assign new_n3692_ = n4545_lo;
  assign new_n3694_ = n4548_lo;
  assign new_n3695_ = ~n4548_lo;
  assign new_n3696_ = n4554_lo;
  assign new_n3698_ = n4557_lo;
  assign new_n3700_ = n4560_lo;
  assign new_n3702_ = n4563_lo;
  assign new_n3703_ = ~n4563_lo;
  assign new_n3704_ = n4566_lo;
  assign new_n3706_ = n4569_lo;
  assign new_n3708_ = n4572_lo;
  assign new_n3710_ = n4575_lo;
  assign new_n3712_ = n4578_lo;
  assign new_n3714_ = n4581_lo;
  assign new_n3716_ = n4584_lo;
  assign new_n3719_ = ~n4587_lo;
  assign new_n3720_ = n4590_lo;
  assign new_n3722_ = n4593_lo;
  assign new_n3724_ = n4596_lo;
  assign new_n3727_ = ~n4599_lo;
  assign new_n3728_ = n4602_lo;
  assign new_n3730_ = n4605_lo;
  assign new_n3732_ = n4608_lo;
  assign new_n3735_ = ~n4611_lo;
  assign new_n3736_ = n4614_lo;
  assign new_n3738_ = n4617_lo;
  assign new_n3740_ = n4620_lo;
  assign new_n3742_ = n4623_lo;
  assign new_n3744_ = n4626_lo;
  assign new_n3746_ = n4629_lo;
  assign new_n3748_ = n4632_lo;
  assign new_n3750_ = n4635_lo;
  assign new_n3752_ = n4638_lo;
  assign new_n3754_ = n4641_lo;
  assign new_n3756_ = n4644_lo;
  assign new_n3758_ = n4647_lo;
  assign new_n3759_ = ~n4647_lo;
  assign new_n3760_ = n4650_lo;
  assign new_n3762_ = n4653_lo;
  assign new_n3764_ = n4656_lo;
  assign new_n3766_ = n4659_lo;
  assign new_n3767_ = ~n4659_lo;
  assign new_n3768_ = n4662_lo;
  assign new_n3770_ = n4665_lo;
  assign new_n3772_ = n4668_lo;
  assign new_n3774_ = n4671_lo;
  assign new_n3775_ = ~n4671_lo;
  assign new_n3776_ = n4674_lo;
  assign new_n3778_ = n4677_lo;
  assign new_n3780_ = n4680_lo;
  assign new_n3782_ = n4683_lo;
  assign new_n3783_ = ~n4683_lo;
  assign new_n3784_ = n4686_lo;
  assign new_n3786_ = n4689_lo;
  assign new_n3788_ = n4692_lo;
  assign new_n3790_ = n4695_lo;
  assign new_n3791_ = ~n4695_lo;
  assign new_n3792_ = n4698_lo;
  assign new_n3794_ = n4701_lo;
  assign new_n3796_ = n4704_lo;
  assign new_n3798_ = n4707_lo;
  assign new_n3799_ = ~n4707_lo;
  assign new_n3800_ = n4710_lo;
  assign new_n3802_ = n4713_lo;
  assign new_n3804_ = n4716_lo;
  assign new_n3806_ = n4719_lo;
  assign new_n3807_ = ~n4719_lo;
  assign new_n3808_ = n4722_lo;
  assign new_n3810_ = n4725_lo;
  assign new_n3812_ = n4728_lo;
  assign new_n3814_ = n4731_lo;
  assign new_n3815_ = ~n4731_lo;
  assign new_n3816_ = n4734_lo;
  assign new_n3818_ = n4737_lo;
  assign new_n3820_ = n4740_lo;
  assign new_n3823_ = ~n4743_lo;
  assign new_n3825_ = ~n6382_o2;
  assign new_n3827_ = ~n6383_o2;
  assign new_n3829_ = ~n6419_o2;
  assign new_n3831_ = ~n6420_o2;
  assign new_n3833_ = ~n6435_o2;
  assign new_n3835_ = ~n6436_o2;
  assign new_n3837_ = ~n6448_o2;
  assign new_n3839_ = ~n6449_o2;
  assign new_n3841_ = ~n6613_o2;
  assign new_n3842_ = n6614_o2;
  assign new_n3845_ = ~n6641_o2;
  assign new_n3846_ = n6658_o2;
  assign new_n3848_ = n6757_o2;
  assign new_n3849_ = ~n6757_o2;
  assign new_n3850_ = n6756_o2;
  assign new_n3851_ = ~n6756_o2;
  assign new_n3853_ = ~n7116_o2;
  assign new_n3854_ = n7156_o2;
  assign new_n3855_ = ~n7156_o2;
  assign new_n3857_ = ~n6549_o2;
  assign new_n3858_ = n6550_o2;
  assign new_n3859_ = ~n6550_o2;
  assign new_n3860_ = n7357_o2;
  assign new_n3862_ = n7358_o2;
  assign new_n3864_ = n7359_o2;
  assign new_n3866_ = n7360_o2;
  assign new_n3868_ = n6621_o2;
  assign new_n3869_ = ~n6621_o2;
  assign new_n3870_ = n6623_o2;
  assign new_n3871_ = ~n6623_o2;
  assign new_n3872_ = n6625_o2;
  assign new_n3873_ = ~n6625_o2;
  assign new_n3874_ = n6626_o2;
  assign new_n3876_ = n6627_o2;
  assign new_n3877_ = ~n6627_o2;
  assign new_n3878_ = n6628_o2;
  assign new_n3880_ = n6629_o2;
  assign new_n3882_ = n6630_o2;
  assign new_n3883_ = ~n6630_o2;
  assign new_n3884_ = n6669_o2;
  assign new_n3885_ = ~n6669_o2;
  assign new_n3886_ = n7449_o2;
  assign new_n3887_ = ~n7449_o2;
  assign new_n3889_ = ~n7450_o2;
  assign new_n3891_ = ~n7451_o2;
  assign new_n3892_ = n7452_o2;
  assign new_n3893_ = ~n7452_o2;
  assign new_n3894_ = n6682_o2;
  assign new_n3895_ = ~n6682_o2;
  assign new_n3896_ = n6683_o2;
  assign new_n3897_ = ~n6683_o2;
  assign new_n3898_ = n6684_o2;
  assign new_n3899_ = ~n6684_o2;
  assign new_n3900_ = n6685_o2;
  assign new_n3901_ = ~n6685_o2;
  assign new_n3902_ = n7463_o2;
  assign new_n3903_ = ~n7463_o2;
  assign new_n3904_ = n6686_o2;
  assign new_n3905_ = ~n6686_o2;
  assign new_n3906_ = n6687_o2;
  assign new_n3907_ = ~n6687_o2;
  assign new_n3908_ = n6688_o2;
  assign new_n3909_ = ~n6688_o2;
  assign new_n3910_ = n6689_o2;
  assign new_n3911_ = ~n6689_o2;
  assign new_n3912_ = n6772_o2;
  assign new_n3913_ = ~n6772_o2;
  assign new_n3914_ = n6773_o2;
  assign new_n3916_ = n6774_o2;
  assign new_n3917_ = ~n6774_o2;
  assign new_n3918_ = n6775_o2;
  assign new_n3919_ = ~n6775_o2;
  assign new_n3921_ = ~G3467_o2;
  assign new_n3922_ = G2810_o2;
  assign new_n3924_ = n6833_o2;
  assign new_n3926_ = n6945_o2;
  assign new_n3927_ = ~n6945_o2;
  assign new_n3928_ = n6947_o2;
  assign new_n3929_ = ~n6947_o2;
  assign new_n3930_ = n6949_o2;
  assign new_n3931_ = ~n6949_o2;
  assign new_n3932_ = n6951_o2;
  assign new_n3934_ = n6888_o2;
  assign new_n3935_ = ~n6888_o2;
  assign new_n3936_ = n6889_o2;
  assign new_n3937_ = ~n6889_o2;
  assign new_n3938_ = n6936_o2;
  assign new_n3939_ = ~n6936_o2;
  assign new_n3940_ = n6954_o2;
  assign new_n3941_ = ~n6954_o2;
  assign new_n3942_ = n6955_o2;
  assign new_n3943_ = ~n6955_o2;
  assign new_n3944_ = n6956_o2;
  assign new_n3945_ = ~n6956_o2;
  assign new_n3946_ = n6957_o2;
  assign new_n3947_ = ~n6957_o2;
  assign new_n3948_ = n6958_o2;
  assign new_n3949_ = ~n6958_o2;
  assign new_n3950_ = n6982_o2;
  assign new_n3951_ = ~n6982_o2;
  assign new_n3952_ = n6984_o2;
  assign new_n3953_ = ~n6984_o2;
  assign new_n3954_ = n6974_o2;
  assign new_n3955_ = ~n6974_o2;
  assign new_n3956_ = n6975_o2;
  assign new_n3957_ = ~n6975_o2;
  assign new_n3958_ = n6999_o2;
  assign new_n3959_ = ~n6999_o2;
  assign new_n3960_ = n7015_o2;
  assign new_n3961_ = ~n7015_o2;
  assign new_n3962_ = n7016_o2;
  assign new_n3963_ = ~n7016_o2;
  assign new_n3964_ = n7017_o2;
  assign new_n3965_ = ~n7017_o2;
  assign new_n3966_ = n7018_o2;
  assign new_n3967_ = ~n7018_o2;
  assign new_n3968_ = n7005_o2;
  assign new_n3969_ = ~n7005_o2;
  assign new_n3970_ = n7019_o2;
  assign new_n3971_ = ~n7019_o2;
  assign new_n3972_ = n7022_o2;
  assign new_n3973_ = ~n7022_o2;
  assign new_n3974_ = n7023_o2;
  assign new_n3975_ = ~n7023_o2;
  assign new_n3976_ = n7132_o2;
  assign new_n3977_ = ~n7132_o2;
  assign new_n3978_ = n7133_o2;
  assign new_n3979_ = ~n7133_o2;
  assign new_n3980_ = n7135_o2;
  assign new_n3981_ = ~n7135_o2;
  assign new_n3982_ = n7136_o2;
  assign new_n3983_ = ~n7136_o2;
  assign new_n3984_ = n7175_o2;
  assign new_n3985_ = ~n7175_o2;
  assign new_n3986_ = n7155_o2;
  assign new_n3987_ = ~n7155_o2;
  assign new_n3989_ = ~G3060_o2;
  assign new_n3990_ = n7383_o2;
  assign new_n3991_ = ~n7383_o2;
  assign new_n3993_ = ~G3802_o2;
  assign new_n3995_ = ~G3859_o2;
  assign new_n3996_ = n7355_o2;
  assign new_n3998_ = n7356_o2;
  assign new_n4001_ = ~G4054_o2;
  assign new_n4003_ = ~G4068_o2;
  assign new_n4004_ = n7384_o2;
  assign new_n4005_ = ~n7384_o2;
  assign new_n4006_ = n7387_o2;
  assign new_n4007_ = ~n7387_o2;
  assign new_n4008_ = n7388_o2;
  assign new_n4010_ = n7389_o2;
  assign new_n4012_ = n7386_o2;
  assign new_n4013_ = ~n7386_o2;
  assign new_n4014_ = n7453_o2;
  assign new_n4015_ = ~n7453_o2;
  assign new_n4016_ = n7431_o2;
  assign new_n4017_ = ~n7431_o2;
  assign new_n4018_ = n7432_o2;
  assign new_n4020_ = n7433_o2;
  assign new_n4022_ = n7430_o2;
  assign new_n4023_ = ~n7430_o2;
  assign new_n4024_ = n7485_o2;
  assign new_n4026_ = n7486_o2;
  assign new_n4028_ = G2508_o2;
  assign new_n4030_ = G2486_o2;
  assign new_n4031_ = ~G2486_o2;
  assign new_n4032_ = n2326_inv;
  assign new_n4034_ = n2329_inv;
  assign new_n4036_ = n3756_lo_buf_o2;
  assign new_n4037_ = ~n3756_lo_buf_o2;
  assign new_n4038_ = n4056_lo_buf_o2;
  assign new_n4040_ = G3474_o2;
  assign new_n4041_ = ~G3474_o2;
  assign new_n4042_ = n2341_inv;
  assign new_n4043_ = ~n2341_inv;
  assign new_n4044_ = n7396_o2;
  assign new_n4046_ = n7398_o2;
  assign new_n4048_ = n7400_o2;
  assign new_n4050_ = n7401_o2;
  assign new_n4052_ = n7402_o2;
  assign new_n4054_ = n7403_o2;
  assign new_n4056_ = n7404_o2;
  assign new_n4058_ = n7405_o2;
  assign new_n4060_ = G2711_o2;
  assign new_n4062_ = n2371_inv;
  assign new_n4064_ = n7490_o2;
  assign new_n4066_ = n7527_o2;
  assign new_n4068_ = n7528_o2;
  assign new_n4070_ = n7529_o2;
  assign new_n4072_ = n7530_o2;
  assign new_n4074_ = n7523_o2;
  assign new_n4076_ = n7524_o2;
  assign new_n4078_ = n7525_o2;
  assign new_n4080_ = n7526_o2;
  assign new_n4082_ = n4296_lo_buf_o2;
  assign new_n4083_ = ~n4296_lo_buf_o2;
  assign new_n4084_ = n4368_lo_buf_o2;
  assign new_n4085_ = ~n4368_lo_buf_o2;
  assign new_n4086_ = G2466_o2;
  assign new_n4087_ = ~G2466_o2;
  assign new_n4088_ = G2404_o2;
  assign new_n4089_ = ~G2404_o2;
  assign new_n4090_ = n7534_o2;
  assign new_n4092_ = n7535_o2;
  assign new_n4094_ = n7536_o2;
  assign new_n4096_ = n7533_o2;
  assign new_n4098_ = G1060_o2;
  assign new_n4099_ = ~G1060_o2;
  assign new_n4100_ = G963_o2;
  assign new_n4101_ = ~G963_o2;
  assign new_n4102_ = G2448_o2;
  assign new_n4104_ = G2685_o2;
  assign new_n4105_ = ~G2685_o2;
  assign new_n4106_ = G2679_o2;
  assign new_n4107_ = ~G2679_o2;
  assign new_n4108_ = G2774_o2;
  assign new_n4109_ = ~G2774_o2;
  assign new_n4110_ = G2780_o2;
  assign new_n4111_ = ~G2780_o2;
  assign new_n4112_ = G2759_o2;
  assign new_n4113_ = ~G2759_o2;
  assign new_n4114_ = G2737_o2;
  assign new_n4116_ = G2850_o2;
  assign new_n4118_ = G3393_o2;
  assign new_n4119_ = ~G3393_o2;
  assign new_n4120_ = G3404_o2;
  assign new_n4121_ = ~G3404_o2;
  assign new_n4122_ = G3559_o2;
  assign new_n4123_ = ~G3559_o2;
  assign new_n4124_ = G2744_o2;
  assign new_n4126_ = n3708_lo_buf_o2;
  assign new_n4128_ = n3840_lo_buf_o2;
  assign new_n4129_ = ~n3840_lo_buf_o2;
  assign new_n4130_ = n4008_lo_buf_o2;
  assign new_n4132_ = n4104_lo_buf_o2;
  assign new_n4134_ = G1821_o2;
  assign new_n4135_ = ~G1821_o2;
  assign new_n4136_ = G1734_o2;
  assign new_n4137_ = ~G1734_o2;
  assign new_n4138_ = G3517_o2;
  assign new_n4140_ = G3533_o2;
  assign new_n4141_ = ~G3533_o2;
  assign new_n4142_ = G3629_o2;
  assign new_n4144_ = G3645_o2;
  assign new_n4145_ = ~G3645_o2;
  assign new_n4146_ = n2497_inv;
  assign new_n4148_ = G2731_o2;
  assign new_n4150_ = G2844_o2;
  assign new_n4152_ = n3732_lo_buf_o2;
  assign new_n4154_ = n4032_lo_buf_o2;
  assign new_n4156_ = G3552_o2;
  assign new_n4157_ = ~G3552_o2;
  assign new_n4158_ = G2271_o2;
  assign new_n4160_ = n4248_lo_buf_o2;
  assign new_n4162_ = n4332_lo_buf_o2;
  assign new_n4164_ = n4344_lo_buf_o2;
  assign new_n4166_ = n4380_lo_buf_o2;
  assign new_n4168_ = G2398_o2;
  assign new_n4170_ = G2480_o2;
  assign new_n4172_ = G2418_o2;
  assign new_n4174_ = G1455_o2;
  assign new_n4175_ = ~G1455_o2;
  assign new_n4176_ = G1449_o2;
  assign new_n4177_ = ~G1449_o2;
  assign new_n4178_ = G1452_o2;
  assign new_n4179_ = ~G1452_o2;
  assign new_n4180_ = G1425_o2;
  assign new_n4181_ = ~G1425_o2;
  assign new_n4182_ = G1428_o2;
  assign new_n4183_ = ~G1428_o2;
  assign new_n4184_ = G1419_o2;
  assign new_n4185_ = ~G1419_o2;
  assign new_n4186_ = G1422_o2;
  assign new_n4187_ = ~G1422_o2;
  assign new_n4188_ = n4308_lo_buf_o2;
  assign new_n4189_ = ~n4308_lo_buf_o2;
  assign new_n4190_ = G2675_o2;
  assign new_n4191_ = ~G2675_o2;
  assign new_n4192_ = G3035_o2;
  assign new_n4193_ = ~G3035_o2;
  assign new_n4194_ = G3026_o2;
  assign new_n4195_ = ~G3026_o2;
  assign new_n4196_ = G3029_o2;
  assign new_n4197_ = ~G3029_o2;
  assign new_n4198_ = G3032_o2;
  assign new_n4199_ = ~G3032_o2;
  assign new_n4200_ = G2999_o2;
  assign new_n4201_ = ~G2999_o2;
  assign new_n4202_ = G3002_o2;
  assign new_n4203_ = ~G3002_o2;
  assign new_n4204_ = G2770_o2;
  assign new_n4205_ = ~G2770_o2;
  assign new_n4206_ = G3008_o2;
  assign new_n4207_ = ~G3008_o2;
  assign new_n4208_ = G2073_o2;
  assign new_n4209_ = ~G2073_o2;
  assign new_n4210_ = G2752_o2;
  assign new_n4211_ = ~G2752_o2;
  assign new_n4212_ = G3005_o2;
  assign new_n4213_ = ~G3005_o2;
  assign new_n4214_ = G5108_o2;
  assign new_n4217_ = ~G5135_o2;
  assign new_n4219_ = ~G5111_o2;
  assign new_n4221_ = ~G5138_o2;
  assign new_n4222_ = G3415_o2;
  assign new_n4223_ = ~G3415_o2;
  assign new_n4224_ = G3386_o2;
  assign new_n4225_ = ~G3386_o2;
  assign new_n4226_ = G3570_o2;
  assign new_n4227_ = ~G3570_o2;
  assign new_n4228_ = G2430_o2;
  assign new_n4229_ = ~G2430_o2;
  assign new_n4230_ = G3495_o2;
  assign new_n4231_ = ~G3495_o2;
  assign new_n4232_ = G3621_o2;
  assign new_n4233_ = ~G3621_o2;
  assign new_n4234_ = n4284_lo_buf_o2;
  assign new_n4235_ = ~n4284_lo_buf_o2;
  assign new_n4236_ = n4356_lo_buf_o2;
  assign new_n4237_ = ~n4356_lo_buf_o2;
  assign new_n4238_ = G2472_o2;
  assign new_n4239_ = ~G2472_o2;
  assign new_n4240_ = G2410_o2;
  assign new_n4241_ = ~G2410_o2;
  assign new_n4242_ = n3960_lo_buf_o2;
  assign new_n4243_ = ~n3960_lo_buf_o2;
  assign new_n4244_ = n3972_lo_buf_o2;
  assign new_n4246_ = n2647_inv;
  assign new_n4247_ = ~n2647_inv;
  assign new_n4248_ = n2650_inv;
  assign new_n4250_ = n3684_lo_buf_o2;
  assign new_n4252_ = n4080_lo_buf_o2;
  assign new_n4253_ = ~n4080_lo_buf_o2;
  assign new_n4254_ = n4092_lo_buf_o2;
  assign new_n4255_ = ~n4092_lo_buf_o2;
  assign new_n4256_ = n2662_inv;
  assign new_n4257_ = ~n2662_inv;
  assign new_n4258_ = n2665_inv;
  assign new_n4259_ = ~n2665_inv;
  assign new_n4260_ = G1147_o2;
  assign new_n4261_ = ~G1147_o2;
  assign new_n4262_ = G2705_o2;
  assign new_n4263_ = ~G2705_o2;
  assign new_n4264_ = G2693_o2;
  assign new_n4265_ = ~G2693_o2;
  assign new_n4266_ = G2696_o2;
  assign new_n4267_ = ~G2696_o2;
  assign new_n4268_ = G2700_o2;
  assign new_n4269_ = ~G2700_o2;
  assign new_n4270_ = G2915_o2;
  assign new_n4271_ = ~G2915_o2;
  assign new_n4272_ = G2966_o2;
  assign new_n4273_ = ~G2966_o2;
  assign new_n4274_ = G2540_o2;
  assign new_n4275_ = ~G2540_o2;
  assign new_n4276_ = G2788_o2;
  assign new_n4277_ = ~G2788_o2;
  assign new_n4278_ = G2792_o2;
  assign new_n4279_ = ~G2792_o2;
  assign new_n4280_ = G2797_o2;
  assign new_n4281_ = ~G2797_o2;
  assign new_n4282_ = G2804_o2;
  assign new_n4283_ = ~G2804_o2;
  assign new_n4284_ = G1038_o2;
  assign new_n4285_ = ~G1038_o2;
  assign new_n4286_ = G1044_o2;
  assign new_n4287_ = ~G1044_o2;
  assign new_n4288_ = G1090_o2;
  assign new_n4289_ = ~G1090_o2;
  assign new_n4290_ = G1096_o2;
  assign new_n4291_ = ~G1096_o2;
  assign new_n4292_ = G1029_o2;
  assign new_n4293_ = ~G1029_o2;
  assign new_n4294_ = G3942_o2;
  assign new_n4295_ = ~G3942_o2;
  assign new_n4296_ = G3954_o2;
  assign new_n4297_ = ~G3954_o2;
  assign new_n4298_ = G4011_o2;
  assign new_n4299_ = ~G4011_o2;
  assign new_n4300_ = G4017_o2;
  assign new_n4301_ = ~G4017_o2;
  assign new_n4302_ = G1141_o2;
  assign new_n4303_ = ~G1141_o2;
  assign new_n4304_ = G1081_o2;
  assign new_n4305_ = ~G1081_o2;
  assign new_n4306_ = G2146_o2;
  assign new_n4307_ = ~G2146_o2;
  assign new_n4308_ = G2145_o2;
  assign new_n4309_ = ~G2145_o2;
  assign new_n4310_ = G2144_o2;
  assign new_n4311_ = ~G2144_o2;
  assign new_n4312_ = G2143_o2;
  assign new_n4313_ = ~G2143_o2;
  assign new_n4314_ = G2142_o2;
  assign new_n4315_ = ~G2142_o2;
  assign new_n4316_ = G2141_o2;
  assign new_n4317_ = ~G2141_o2;
  assign new_n4318_ = G2140_o2;
  assign new_n4319_ = ~G2140_o2;
  assign new_n4320_ = G2139_o2;
  assign new_n4321_ = ~G2139_o2;
  assign new_n4322_ = G3769_o2;
  assign new_n4323_ = ~G3769_o2;
  assign new_n4324_ = G3773_o2;
  assign new_n4325_ = ~G3773_o2;
  assign new_n4326_ = G3768_o2;
  assign new_n4327_ = ~G3768_o2;
  assign new_n4328_ = G4101_o2;
  assign new_n4329_ = ~G4101_o2;
  assign new_n4330_ = G3161_o2;
  assign new_n4331_ = ~G3161_o2;
  assign new_n4332_ = G4143_o2;
  assign new_n4333_ = ~G4143_o2;
  assign new_n4334_ = G3828_o2;
  assign new_n4335_ = ~G3828_o2;
  assign new_n4336_ = G3831_o2;
  assign new_n4337_ = ~G3831_o2;
  assign new_n4338_ = G3334_o2;
  assign new_n4339_ = ~G3334_o2;
  assign new_n4340_ = G3335_o2;
  assign new_n4341_ = ~G3335_o2;
  assign new_n4342_ = G3180_o2;
  assign new_n4343_ = ~G3180_o2;
  assign new_n4344_ = G3340_o2;
  assign new_n4345_ = ~G3340_o2;
  assign new_n4346_ = G3339_o2;
  assign new_n4347_ = ~G3339_o2;
  assign new_n4348_ = G3341_o2;
  assign new_n4349_ = ~G3341_o2;
  assign new_n4350_ = G3234_o2;
  assign new_n4351_ = ~G3234_o2;
  assign new_n4352_ = G3829_o2;
  assign new_n4353_ = ~G3829_o2;
  assign new_n4354_ = G3338_o2;
  assign new_n4355_ = ~G3338_o2;
  assign new_n4356_ = G3336_o2;
  assign new_n4357_ = ~G3336_o2;
  assign new_n4358_ = G3770_o2;
  assign new_n4359_ = ~G3770_o2;
  assign new_n4360_ = G3918_o2;
  assign new_n4361_ = ~G3918_o2;
  assign new_n4362_ = G3774_o2;
  assign new_n4363_ = ~G3774_o2;
  assign new_n4364_ = G3921_o2;
  assign new_n4365_ = ~G3921_o2;
  assign new_n4366_ = G3832_o2;
  assign new_n4367_ = ~G3832_o2;
  assign new_n4368_ = G3993_o2;
  assign new_n4369_ = ~G3993_o2;
  assign new_n4370_ = G2076_o2;
  assign new_n4371_ = ~G2076_o2;
  assign new_n4372_ = G2071_o2;
  assign new_n4373_ = ~G2071_o2;
  assign new_n4374_ = G2072_o2;
  assign new_n4375_ = ~G2072_o2;
  assign new_n4376_ = G2069_o2;
  assign new_n4377_ = ~G2069_o2;
  assign new_n4378_ = G2070_o2;
  assign new_n4379_ = ~G2070_o2;
  assign new_n4380_ = G2067_o2;
  assign new_n4381_ = ~G2067_o2;
  assign new_n4382_ = G2068_o2;
  assign new_n4383_ = ~G2068_o2;
  assign new_n4384_ = G4095_o2;
  assign new_n4385_ = ~G4095_o2;
  assign new_n4386_ = G3272_o2;
  assign new_n4387_ = ~G3272_o2;
  assign new_n4388_ = G3269_o2;
  assign new_n4389_ = ~G3269_o2;
  assign new_n4390_ = G3270_o2;
  assign new_n4391_ = ~G3270_o2;
  assign new_n4392_ = G3271_o2;
  assign new_n4393_ = ~G3271_o2;
  assign new_n4394_ = G3265_o2;
  assign new_n4395_ = ~G3265_o2;
  assign new_n4396_ = G3266_o2;
  assign new_n4397_ = ~G3266_o2;
  assign new_n4398_ = G4137_o2;
  assign new_n4399_ = ~G4137_o2;
  assign new_n4400_ = G3268_o2;
  assign new_n4401_ = ~G3268_o2;
  assign new_n4402_ = G2361_o2;
  assign new_n4403_ = ~G2361_o2;
  assign new_n4404_ = G3228_o2;
  assign new_n4405_ = ~G3228_o2;
  assign new_n4406_ = G3267_o2;
  assign new_n4407_ = ~G3267_o2;
  assign new_n4408_ = G2336_o2;
  assign new_n4409_ = ~G2336_o2;
  assign new_n4410_ = G3459_o2;
  assign new_n4411_ = ~G3459_o2;
  assign new_n4412_ = G3428_o2;
  assign new_n4413_ = ~G3428_o2;
  assign new_n4414_ = G3438_o2;
  assign new_n4415_ = ~G3438_o2;
  assign new_n4416_ = G3449_o2;
  assign new_n4417_ = ~G3449_o2;
  assign new_n4418_ = G3421_o2;
  assign new_n4419_ = ~G3421_o2;
  assign new_n4420_ = G3576_o2;
  assign new_n4421_ = ~G3576_o2;
  assign new_n4422_ = G3303_o2;
  assign new_n4423_ = ~G3303_o2;
  assign new_n4424_ = G3583_o2;
  assign new_n4425_ = ~G3583_o2;
  assign new_n4426_ = G3594_o2;
  assign new_n4427_ = ~G3594_o2;
  assign new_n4428_ = G3674_o2;
  assign new_n4429_ = ~G3674_o2;
  assign new_n4430_ = G3685_o2;
  assign new_n4431_ = ~G3685_o2;
  assign new_n4432_ = G4504_o2;
  assign new_n4433_ = ~G4504_o2;
  assign new_n4434_ = G4180_o2;
  assign new_n4435_ = ~G4180_o2;
  assign new_n4437_ = ~G5123_o2;
  assign new_n4438_ = G5142_o2;
  assign new_n4440_ = G5126_o2;
  assign new_n4442_ = G5144_o2;
  assign new_n4444_ = G3912_o2;
  assign new_n4445_ = ~G3912_o2;
  assign new_n4446_ = G4417_o2;
  assign new_n4447_ = ~G4417_o2;
  assign new_n4448_ = G4420_o2;
  assign new_n4449_ = ~G4420_o2;
  assign new_n4450_ = G3969_o2;
  assign new_n4451_ = ~G3969_o2;
  assign new_n4452_ = G4023_o2;
  assign new_n4453_ = ~G4023_o2;
  assign new_n4454_ = G2720_o2;
  assign new_n4455_ = ~G2720_o2;
  assign new_n4456_ = G2837_o2;
  assign new_n4457_ = ~G2837_o2;
  assign new_n4458_ = n2965_inv;
  assign new_n4459_ = ~n2965_inv;
  assign new_n4460_ = n2968_inv;
  assign new_n4461_ = ~n2968_inv;
  assign new_n4462_ = n2971_inv;
  assign new_n4463_ = ~n2971_inv;
  assign new_n4464_ = n2974_inv;
  assign new_n4465_ = ~n2974_inv;
  assign new_n4466_ = G1876_o2;
  assign new_n4467_ = ~G1876_o2;
  assign new_n4468_ = G4996_o2;
  assign new_n4469_ = ~G4996_o2;
  assign new_n4470_ = G4984_o2;
  assign new_n4471_ = ~G4984_o2;
  assign new_n4472_ = G4920_o2;
  assign new_n4473_ = ~G4920_o2;
  assign new_n4474_ = G4923_o2;
  assign new_n4475_ = ~G4923_o2;
  assign new_n4476_ = G4930_o2;
  assign new_n4477_ = ~G4930_o2;
  assign new_n4478_ = G4933_o2;
  assign new_n4479_ = ~G4933_o2;
  assign new_n4480_ = n4320_lo_buf_o2;
  assign new_n4481_ = ~n4320_lo_buf_o2;
  assign new_n4482_ = G2424_o2;
  assign new_n4483_ = ~G2424_o2;
  assign new_n4484_ = G3317_o2;
  assign new_n4486_ = G3503_o2;
  assign new_n4488_ = G3485_o2;
  assign new_n4489_ = ~G3485_o2;
  assign new_n4490_ = G3611_o2;
  assign new_n4491_ = ~G3611_o2;
  assign new_n4492_ = n3864_lo_buf_o2;
  assign new_n4494_ = n3888_lo_buf_o2;
  assign new_n4496_ = n4116_lo_buf_o2;
  assign new_n4498_ = n4128_lo_buf_o2;
  assign new_n4500_ = n4140_lo_buf_o2;
  assign new_n4502_ = n4152_lo_buf_o2;
  assign new_n4504_ = G1815_o2;
  assign new_n4505_ = ~G1815_o2;
  assign new_n4506_ = G1728_o2;
  assign new_n4507_ = ~G1728_o2;
  assign new_n4508_ = G1035_o2;
  assign new_n4509_ = ~G1035_o2;
  assign new_n4510_ = G1041_o2;
  assign new_n4511_ = ~G1041_o2;
  assign new_n4512_ = G1087_o2;
  assign new_n4513_ = ~G1087_o2;
  assign new_n4514_ = G1093_o2;
  assign new_n4515_ = ~G1093_o2;
  assign new_n4516_ = G1132_o2;
  assign new_n4517_ = ~G1132_o2;
  assign new_n4518_ = G1108_o2;
  assign new_n4519_ = ~G1108_o2;
  assign new_n4520_ = G1138_o2;
  assign new_n4521_ = ~G1138_o2;
  assign new_n4522_ = G1114_o2;
  assign new_n4523_ = ~G1114_o2;
  assign new_n4524_ = G1807_o2;
  assign new_n4525_ = ~G1807_o2;
  assign new_n4526_ = G2108_o2;
  assign new_n4527_ = ~G2108_o2;
  assign new_n4528_ = G1126_o2;
  assign new_n4529_ = ~G1126_o2;
  assign new_n4530_ = G1899_o2;
  assign new_n4531_ = ~G1899_o2;
  assign new_n4532_ = G2134_o2;
  assign new_n4533_ = ~G2134_o2;
  assign new_n4534_ = G1852_o2;
  assign new_n4535_ = ~G1852_o2;
  assign new_n4536_ = G2116_o2;
  assign new_n4537_ = ~G2116_o2;
  assign new_n4538_ = G2543_o2;
  assign new_n4539_ = ~G2543_o2;
  assign new_n4540_ = G2727_o2;
  assign new_n4541_ = ~G2727_o2;
  assign new_n4542_ = G2715_o2;
  assign new_n4543_ = ~G2715_o2;
  assign new_n4544_ = G2832_o2;
  assign new_n4545_ = ~G2832_o2;
  assign new_n4546_ = G1873_o2;
  assign new_n4547_ = ~G1873_o2;
  assign new_n4548_ = G3291_o2;
  assign new_n4549_ = ~G3291_o2;
  assign new_n4550_ = G5025_o2;
  assign new_n4551_ = ~G5025_o2;
  assign new_n4552_ = G5036_o2;
  assign new_n4553_ = ~G5036_o2;
  assign new_n4554_ = G3132_o2;
  assign new_n4555_ = ~G3132_o2;
  assign new_n4556_ = G5038_o2;
  assign new_n4557_ = ~G5038_o2;
  assign new_n4558_ = G5039_o2;
  assign new_n4559_ = ~G5039_o2;
  assign new_n4560_ = n3118_inv;
  assign new_n4561_ = ~n3118_inv;
  assign new_n4562_ = n3121_inv;
  assign new_n4563_ = ~n3121_inv;
  assign new_n4564_ = n3124_inv;
  assign new_n4565_ = ~n3124_inv;
  assign new_n4566_ = n3127_inv;
  assign new_n4567_ = ~n3127_inv;
  assign new_n4568_ = n3984_lo_buf_o2;
  assign new_n4570_ = G1802_o2;
  assign new_n4571_ = ~G1802_o2;
  assign new_n4572_ = G1804_o2;
  assign new_n4573_ = ~G1804_o2;
  assign new_n4574_ = G1849_o2;
  assign new_n4575_ = ~G1849_o2;
  assign new_n4576_ = G1851_o2;
  assign new_n4577_ = ~G1851_o2;
  assign new_n4578_ = G2492_o2;
  assign new_n4579_ = ~G2492_o2;
  assign new_n4580_ = G1799_o2;
  assign new_n4581_ = ~G1799_o2;
  assign new_n4582_ = G4231_o2;
  assign new_n4583_ = ~G4231_o2;
  assign new_n4584_ = G4234_o2;
  assign new_n4585_ = ~G4234_o2;
  assign new_n4586_ = G4245_o2;
  assign new_n4587_ = ~G4245_o2;
  assign new_n4588_ = G4247_o2;
  assign new_n4589_ = ~G4247_o2;
  assign new_n4590_ = G1894_o2;
  assign new_n4591_ = ~G1894_o2;
  assign new_n4592_ = G1846_o2;
  assign new_n4593_ = ~G1846_o2;
  assign new_n4594_ = G4238_o2;
  assign new_n4595_ = ~G4238_o2;
  assign new_n4596_ = G4249_o2;
  assign new_n4597_ = ~G4249_o2;
  assign new_n4598_ = G2293_o2;
  assign new_n4599_ = ~G2293_o2;
  assign new_n4600_ = G5022_o2;
  assign new_n4601_ = ~G5022_o2;
  assign new_n4602_ = G5006_o2;
  assign new_n4603_ = ~G5006_o2;
  assign new_n4604_ = G4944_o2;
  assign new_n4605_ = ~G4944_o2;
  assign new_n4606_ = G4946_o2;
  assign new_n4607_ = ~G4946_o2;
  assign new_n4608_ = G4954_o2;
  assign new_n4609_ = ~G4954_o2;
  assign new_n4610_ = G4956_o2;
  assign new_n4611_ = ~G4956_o2;
  assign new_n4612_ = G3546_o2;
  assign new_n4613_ = ~G3546_o2;
  assign new_n4614_ = G3658_o2;
  assign new_n4615_ = ~G3658_o2;
  assign new_n4616_ = G1344_o2;
  assign new_n4617_ = ~G1344_o2;
  assign new_n4618_ = G2921_o2;
  assign new_n4619_ = ~G2921_o2;
  assign new_n4620_ = n3912_lo_buf_o2;
  assign new_n4622_ = G1835_o2;
  assign new_n4623_ = ~G1835_o2;
  assign new_n4624_ = G3810_o2;
  assign new_n4625_ = ~G3810_o2;
  assign new_n4626_ = G3866_o2;
  assign new_n4627_ = ~G3866_o2;
  assign new_n4628_ = G3811_o2;
  assign new_n4629_ = ~G3811_o2;
  assign new_n4630_ = G2269_o2;
  assign new_n4631_ = ~G2269_o2;
  assign new_n4632_ = G3812_o2;
  assign new_n4633_ = ~G3812_o2;
  assign new_n4634_ = G3867_o2;
  assign new_n4635_ = ~G3867_o2;
  assign new_n4636_ = G3868_o2;
  assign new_n4637_ = ~G3868_o2;
  assign new_n4638_ = G3809_o2;
  assign new_n4639_ = ~G3809_o2;
  assign new_n4640_ = G3716_o2;
  assign new_n4641_ = ~G3716_o2;
  assign new_n4642_ = G4529_o2;
  assign new_n4643_ = ~G4529_o2;
  assign new_n4644_ = G4670_o2;
  assign new_n4645_ = ~G4670_o2;
  assign new_n4646_ = G4493_o2;
  assign new_n4647_ = ~G4493_o2;
  assign new_n4648_ = G4580_o2;
  assign new_n4649_ = ~G4580_o2;
  assign new_n4650_ = G3822_o2;
  assign new_n4651_ = ~G3822_o2;
  assign new_n4652_ = G3877_o2;
  assign new_n4653_ = ~G3877_o2;
  assign new_n4654_ = G4131_o2;
  assign new_n4655_ = ~G4131_o2;
  assign new_n4656_ = G4170_o2;
  assign new_n4657_ = ~G4170_o2;
  assign new_n4658_ = G4051_o2;
  assign new_n4659_ = ~G4051_o2;
  assign new_n4660_ = G4065_o2;
  assign new_n4661_ = ~G4065_o2;
  assign new_n4662_ = G4697_o2;
  assign new_n4663_ = ~G4697_o2;
  assign new_n4664_ = G4706_o2;
  assign new_n4665_ = ~G4706_o2;
  assign new_n4666_ = G2460_o2;
  assign new_n4667_ = ~G2460_o2;
  assign new_n4668_ = G2454_o2;
  assign new_n4669_ = ~G2454_o2;
  assign new_n4670_ = G2392_o2;
  assign new_n4671_ = ~G2392_o2;
  assign new_n4672_ = G2386_o2;
  assign new_n4673_ = ~G2386_o2;
  assign new_n4674_ = n4260_lo_buf_o2;
  assign new_n4675_ = ~n4260_lo_buf_o2;
  assign new_n4676_ = n4272_lo_buf_o2;
  assign new_n4677_ = ~n4272_lo_buf_o2;
  assign new_n4678_ = n4392_lo_buf_o2;
  assign new_n4679_ = ~n4392_lo_buf_o2;
  assign new_n4680_ = n4404_lo_buf_o2;
  assign new_n4681_ = ~n4404_lo_buf_o2;
  assign new_n4682_ = G1512_o2;
  assign new_n4683_ = ~G1512_o2;
  assign new_n4684_ = G3135_o2;
  assign new_n4685_ = ~G3135_o2;
  assign new_n4686_ = G2379_o2;
  assign new_n4687_ = ~G2379_o2;
  assign new_n4688_ = n4164_lo_buf_o2;
  assign new_n4689_ = ~n4164_lo_buf_o2;
  assign new_n4690_ = n4176_lo_buf_o2;
  assign new_n4691_ = ~n4176_lo_buf_o2;
  assign new_n4692_ = n4224_lo_buf_o2;
  assign new_n4693_ = ~n4224_lo_buf_o2;
  assign new_n4694_ = G2975_o2;
  assign new_n4695_ = ~G2975_o2;
  assign new_n4696_ = G2978_o2;
  assign new_n4697_ = ~G2978_o2;
  assign new_n4698_ = G2933_o2;
  assign new_n4699_ = ~G2933_o2;
  assign new_n4700_ = G2936_o2;
  assign new_n4701_ = ~G2936_o2;
  assign new_n4702_ = G1356_o2;
  assign new_n4703_ = ~G1356_o2;
  assign new_n4704_ = G1359_o2;
  assign new_n4705_ = ~G1359_o2;
  assign new_n4706_ = G1398_o2;
  assign new_n4707_ = ~G1398_o2;
  assign new_n4708_ = G1401_o2;
  assign new_n4709_ = ~G1401_o2;
  assign new_n4710_ = new_n3650_ & new_n3626_;
  assign new_n4711_ = new_n3218_ & new_n8443_;
  assign new_n4712_ = new_n3538_ & new_n8444_;
  assign new_n4713_ = new_n8445_ & new_n3186_;
  assign new_n4714_ = new_n3710_ | new_n8446_;
  assign new_n4715_ = new_n8447_ | new_n8448_;
  assign new_n4716_ = new_n2778_ & new_n2770_;
  assign new_n4717_ = new_n2779_ | new_n8446_;
  assign new_n4718_ = new_n8452_ | new_n3203_;
  assign new_n4719_ = new_n8463_ | new_n2955_;
  assign new_n4720_ = new_n8470_ | new_n2947_;
  assign new_n4721_ = new_n4720_ & new_n4719_;
  assign new_n4722_ = new_n4721_ | new_n8452_;
  assign new_n4723_ = new_n8463_ | new_n2787_;
  assign new_n4724_ = new_n8470_ | new_n2963_;
  assign new_n4725_ = new_n4724_ & new_n4723_;
  assign new_n4726_ = new_n4725_ | new_n8453_;
  assign new_n4727_ = new_n8464_ | new_n8475_;
  assign new_n4728_ = new_n8471_ | new_n8475_;
  assign new_n4729_ = new_n4728_ & new_n4727_;
  assign new_n4730_ = new_n4729_ | new_n8453_;
  assign new_n4731_ = new_n8464_ | new_n2747_;
  assign new_n4732_ = new_n4731_ | new_n8455_;
  assign new_n4733_ = new_n8471_ | new_n2755_;
  assign new_n4734_ = new_n4733_ | new_n8455_;
  assign new_n4735_ = new_n8476_ | new_n8466_;
  assign new_n4736_ = new_n8476_ | new_n8473_;
  assign new_n4737_ = new_n4734_ & new_n4732_;
  assign new_n4738_ = new_n4737_ & new_n8478_;
  assign new_n4739_ = new_n4738_ & new_n8481_;
  assign new_n4740_ = new_n4739_ | new_n8485_;
  assign new_n4741_ = new_n8466_ | new_n2763_;
  assign new_n4742_ = new_n4741_ | new_n8456_;
  assign new_n4743_ = new_n8473_ | new_n2923_;
  assign new_n4744_ = new_n4743_ | new_n8456_;
  assign new_n4745_ = new_n4744_ & new_n4742_;
  assign new_n4746_ = new_n4745_ & new_n8478_;
  assign new_n4747_ = new_n4746_ & new_n8481_;
  assign new_n4748_ = new_n4747_ | new_n8485_;
  assign new_n4749_ = new_n8467_ | new_n2907_;
  assign new_n4750_ = new_n4749_ | new_n8459_;
  assign new_n4751_ = new_n8474_ | new_n2739_;
  assign new_n4752_ = new_n4751_ | new_n8459_;
  assign new_n4753_ = new_n4752_ & new_n4750_;
  assign new_n4754_ = new_n4753_ & new_n8479_;
  assign new_n4755_ = new_n4754_ & new_n8482_;
  assign new_n4756_ = new_n4755_ | new_n8484_;
  assign new_n4757_ = new_n8467_ | new_n2931_;
  assign new_n4758_ = new_n4757_ | new_n8458_;
  assign new_n4759_ = new_n8474_ | new_n2915_;
  assign new_n4760_ = new_n4759_ | new_n8460_;
  assign new_n4761_ = new_n4760_ & new_n4758_;
  assign new_n4762_ = new_n4761_ & new_n8479_;
  assign new_n4763_ = new_n4762_ & new_n8482_;
  assign new_n4764_ = new_n4763_ | new_n8486_;
  assign new_n4765_ = new_n8488_ | new_n8489_;
  assign new_n4766_ = new_n4765_ | new_n8490_;
  assign new_n4767_ = new_n8492_ | new_n8489_;
  assign new_n4768_ = new_n4767_ | new_n8493_;
  assign new_n4769_ = new_n4768_ & new_n4766_;
  assign new_n4770_ = new_n8495_ & new_n8493_;
  assign new_n4771_ = new_n8497_ & new_n8490_;
  assign new_n4772_ = new_n4771_ | new_n4770_;
  assign new_n4773_ = new_n4772_ | new_n3588_;
  assign new_n4774_ = new_n4773_ & new_n4769_;
  assign new_n4775_ = new_n8488_ | new_n8498_;
  assign new_n4776_ = new_n4775_ | new_n8499_;
  assign new_n4777_ = new_n8492_ | new_n8498_;
  assign new_n4778_ = new_n4777_ | new_n8500_;
  assign new_n4779_ = new_n4778_ & new_n4776_;
  assign new_n4780_ = new_n8495_ & new_n8500_;
  assign new_n4781_ = new_n8497_ & new_n8499_;
  assign new_n4782_ = new_n4781_ | new_n4780_;
  assign new_n4783_ = new_n4782_ | new_n3584_;
  assign new_n4784_ = new_n4783_ & new_n4779_;
  assign new_n4785_ = new_n8487_ | new_n3478_;
  assign new_n4786_ = new_n8491_ | new_n3479_;
  assign new_n4787_ = new_n4786_ & new_n4785_;
  assign new_n4788_ = new_n8494_ & new_n8502_;
  assign new_n4789_ = new_n3886_ | new_n8503_;
  assign new_n4790_ = new_n8496_ & new_n8503_;
  assign new_n4791_ = new_n3892_ | new_n8502_;
  assign new_n4792_ = new_n4791_ & new_n4789_;
  assign new_n4793_ = new_n4790_ | new_n4788_;
  assign new_n4794_ = new_n8504_ | new_n8505_;
  assign new_n4795_ = new_n4794_ | new_n8506_;
  assign new_n4796_ = new_n4795_ | new_n4793_;
  assign new_n4797_ = new_n8510_ | new_n8518_;
  assign new_n4798_ = new_n4797_ | new_n8519_;
  assign new_n4799_ = new_n8523_ | new_n8518_;
  assign new_n4800_ = new_n4799_ | new_n8530_;
  assign new_n4801_ = new_n4800_ & new_n4798_;
  assign new_n4802_ = new_n8534_ & new_n8530_;
  assign new_n4803_ = new_n8545_ & new_n8519_;
  assign new_n4804_ = new_n4803_ | new_n4802_;
  assign new_n4805_ = new_n4804_ | new_n3602_;
  assign new_n4806_ = new_n4805_ & new_n4801_;
  assign new_n4807_ = new_n8510_ | new_n8552_;
  assign new_n4808_ = new_n4807_ | new_n8553_;
  assign new_n4809_ = new_n8523_ | new_n8552_;
  assign new_n4810_ = new_n4809_ | new_n8554_;
  assign new_n4811_ = new_n4810_ & new_n4808_;
  assign new_n4812_ = new_n8534_ & new_n8554_;
  assign new_n4813_ = new_n8545_ & new_n8553_;
  assign new_n4814_ = new_n4813_ | new_n4812_;
  assign new_n4815_ = new_n4814_ | new_n3600_;
  assign new_n4816_ = new_n4815_ & new_n4811_;
  assign new_n4817_ = new_n8511_ | new_n3599_;
  assign new_n4818_ = new_n8535_ | new_n3598_;
  assign new_n4819_ = new_n4818_ & new_n4817_;
  assign new_n4820_ = new_n8511_ | new_n8556_;
  assign new_n4821_ = new_n4820_ | new_n8557_;
  assign new_n4822_ = new_n8524_ | new_n8556_;
  assign new_n4823_ = new_n4822_ | new_n8558_;
  assign new_n4824_ = new_n4823_ & new_n4821_;
  assign new_n4825_ = new_n8535_ & new_n8558_;
  assign new_n4826_ = new_n8546_ & new_n8557_;
  assign new_n4827_ = new_n4826_ | new_n4825_;
  assign new_n4828_ = new_n4827_ | new_n8559_;
  assign new_n4829_ = new_n4828_ & new_n4824_;
  assign new_n4830_ = new_n8560_ | new_n8561_;
  assign new_n4831_ = new_n4830_ | new_n8562_;
  assign new_n4832_ = new_n4831_ | new_n8563_;
  assign new_n4833_ = new_n4832_ | new_n4796_;
  assign new_n4834_ = new_n4833_ | new_n4028_;
  assign new_n4835_ = new_n8513_ | new_n8565_;
  assign new_n4836_ = new_n4835_ | new_n8566_;
  assign new_n4837_ = new_n8524_ | new_n8565_;
  assign new_n4838_ = new_n4837_ | new_n8567_;
  assign new_n4839_ = new_n4838_ & new_n4836_;
  assign new_n4840_ = new_n8537_ & new_n8567_;
  assign new_n4841_ = new_n8546_ & new_n8566_;
  assign new_n4842_ = new_n4841_ | new_n4840_;
  assign new_n4843_ = new_n4842_ | new_n8568_;
  assign new_n4844_ = new_n4843_ & new_n4839_;
  assign new_n4845_ = new_n8513_ | new_n8569_;
  assign new_n4846_ = new_n4845_ | new_n8570_;
  assign new_n4847_ = new_n8526_ | new_n8569_;
  assign new_n4848_ = new_n4847_ | new_n8571_;
  assign new_n4849_ = new_n4848_ & new_n4846_;
  assign new_n4850_ = new_n8537_ & new_n8571_;
  assign new_n4851_ = new_n8548_ & new_n8570_;
  assign new_n4852_ = new_n4851_ | new_n4850_;
  assign new_n4853_ = new_n4852_ | new_n3560_;
  assign new_n4854_ = new_n4853_ & new_n4849_;
  assign new_n4855_ = new_n8514_ | new_n8572_;
  assign new_n4856_ = new_n4855_ | new_n8573_;
  assign new_n4857_ = new_n8526_ | new_n8572_;
  assign new_n4858_ = new_n4857_ | new_n8574_;
  assign new_n4859_ = new_n4858_ & new_n4856_;
  assign new_n4860_ = new_n8538_ & new_n8574_;
  assign new_n4861_ = new_n8548_ & new_n8573_;
  assign new_n4862_ = new_n4861_ | new_n4860_;
  assign new_n4863_ = new_n4862_ | new_n3580_;
  assign new_n4864_ = new_n4863_ & new_n4859_;
  assign new_n4865_ = new_n8514_ | new_n8575_;
  assign new_n4866_ = new_n4865_ | new_n8576_;
  assign new_n4867_ = new_n8525_ | new_n8575_;
  assign new_n4868_ = new_n4867_ | new_n8577_;
  assign new_n4869_ = new_n4868_ & new_n4866_;
  assign new_n4870_ = new_n8538_ & new_n8577_;
  assign new_n4871_ = new_n8547_ & new_n8576_;
  assign new_n4872_ = new_n4871_ | new_n4870_;
  assign new_n4873_ = new_n4872_ | new_n3576_;
  assign new_n4874_ = new_n4873_ & new_n4869_;
  assign new_n4875_ = new_n8578_ | new_n8579_;
  assign new_n4876_ = new_n4875_ | new_n8580_;
  assign new_n4877_ = new_n4876_ | new_n8581_;
  assign new_n4878_ = new_n8516_ | new_n8582_;
  assign new_n4879_ = new_n4878_ | new_n8583_;
  assign new_n4880_ = new_n8528_ | new_n8582_;
  assign new_n4881_ = new_n4880_ | new_n8584_;
  assign new_n4882_ = new_n4881_ & new_n4879_;
  assign new_n4883_ = new_n8540_ & new_n8584_;
  assign new_n4884_ = new_n8550_ & new_n8583_;
  assign new_n4885_ = new_n4884_ | new_n4883_;
  assign new_n4886_ = new_n4885_ | new_n3540_;
  assign new_n4887_ = new_n4886_ & new_n4882_;
  assign new_n4888_ = new_n8516_ | new_n8585_;
  assign new_n4889_ = new_n4888_ | new_n8586_;
  assign new_n4890_ = new_n8528_ | new_n8585_;
  assign new_n4891_ = new_n4890_ | new_n8587_;
  assign new_n4892_ = new_n4891_ & new_n4889_;
  assign new_n4893_ = new_n8540_ & new_n8587_;
  assign new_n4894_ = new_n8550_ & new_n8586_;
  assign new_n4895_ = new_n4894_ | new_n4893_;
  assign new_n4896_ = new_n4895_ | new_n3556_;
  assign new_n4897_ = new_n4896_ & new_n4892_;
  assign new_n4898_ = new_n8517_ | new_n8588_;
  assign new_n4899_ = new_n4898_ | new_n8589_;
  assign new_n4900_ = new_n8529_ | new_n8588_;
  assign new_n4901_ = new_n4900_ | new_n8590_;
  assign new_n4902_ = new_n4901_ & new_n4899_;
  assign new_n4903_ = new_n8541_ & new_n8590_;
  assign new_n4904_ = new_n8551_ & new_n8589_;
  assign new_n4905_ = new_n4904_ | new_n4903_;
  assign new_n4906_ = new_n4905_ | new_n3554_;
  assign new_n4907_ = new_n4906_ & new_n4902_;
  assign new_n4908_ = new_n8517_ | new_n8591_;
  assign new_n4909_ = new_n4908_ | new_n8592_;
  assign new_n4910_ = new_n8529_ | new_n8591_;
  assign new_n4911_ = new_n4910_ | new_n8593_;
  assign new_n4912_ = new_n4911_ & new_n4909_;
  assign new_n4913_ = new_n8541_ & new_n8593_;
  assign new_n4914_ = new_n8551_ & new_n8592_;
  assign new_n4915_ = new_n4914_ | new_n4913_;
  assign new_n4916_ = new_n4915_ | new_n3552_;
  assign new_n4917_ = new_n4916_ & new_n4912_;
  assign new_n4918_ = new_n8594_ | new_n8595_;
  assign new_n4919_ = new_n4918_ | new_n8596_;
  assign new_n4920_ = new_n4919_ | new_n8597_;
  assign new_n4921_ = new_n4920_ | new_n4877_;
  assign new_n4922_ = new_n4921_ | new_n3989_;
  assign new_n4923_ = new_n3837_ | new_n8598_;
  assign new_n4924_ = new_n4923_ | new_n8600_;
  assign new_n4925_ = new_n4924_ | new_n8602_;
  assign new_n4926_ = new_n8604_ | new_n3993_;
  assign new_n4927_ = new_n8605_ | new_n8607_;
  assign new_n4928_ = new_n4927_ | new_n8610_;
  assign new_n4929_ = new_n4928_ | new_n8613_;
  assign new_n4930_ = new_n8619_ & new_n8625_;
  assign new_n4931_ = new_n8629_ | new_n8635_;
  assign new_n4932_ = new_n4930_ & new_n8638_;
  assign new_n4933_ = new_n4931_ | new_n8643_;
  assign new_n4934_ = new_n4932_ & new_n8648_;
  assign new_n4935_ = new_n4933_ | new_n8653_;
  assign new_n4936_ = new_n4934_ & new_n8658_;
  assign new_n4937_ = new_n4935_ | new_n8663_;
  assign new_n4938_ = new_n8666_ | new_n8667_;
  assign new_n4939_ = new_n3839_ | new_n8668_;
  assign new_n4940_ = new_n4939_ | new_n8670_;
  assign new_n4941_ = new_n4940_ | new_n8672_;
  assign new_n4942_ = new_n8674_ | new_n3995_;
  assign new_n4943_ = new_n8675_ | new_n8677_;
  assign new_n4944_ = new_n4943_ | new_n8680_;
  assign new_n4945_ = new_n4944_ | new_n8683_;
  assign new_n4946_ = new_n8688_ & new_n8694_;
  assign new_n4947_ = new_n8698_ | new_n8704_;
  assign new_n4948_ = new_n4946_ & new_n8707_;
  assign new_n4949_ = new_n4947_ | new_n8712_;
  assign new_n4950_ = new_n4948_ & new_n8717_;
  assign new_n4951_ = new_n4949_ | new_n8722_;
  assign new_n4952_ = new_n4950_ & new_n8727_;
  assign new_n4953_ = new_n4951_ | new_n8732_;
  assign new_n4954_ = new_n8735_ | new_n8736_;
  assign new_n4955_ = new_n4380_ & new_n4187_;
  assign new_n4956_ = new_n4381_ | new_n4186_;
  assign new_n4957_ = new_n4382_ & new_n4185_;
  assign new_n4958_ = new_n4383_ | new_n4184_;
  assign new_n4959_ = new_n4958_ & new_n4956_;
  assign new_n4960_ = new_n4957_ | new_n4955_;
  assign new_n4961_ = new_n4376_ & new_n4183_;
  assign new_n4962_ = new_n4377_ | new_n4182_;
  assign new_n4963_ = new_n4378_ & new_n4181_;
  assign new_n4964_ = new_n4379_ | new_n4180_;
  assign new_n4965_ = new_n4964_ & new_n4962_;
  assign new_n4966_ = new_n4963_ | new_n4961_;
  assign new_n4967_ = new_n8737_ & new_n8738_;
  assign new_n4968_ = new_n8739_ | new_n8740_;
  assign new_n4969_ = new_n8739_ & new_n8740_;
  assign new_n4970_ = new_n8737_ | new_n8738_;
  assign new_n4971_ = new_n4970_ & new_n4968_;
  assign new_n4972_ = new_n4969_ | new_n4967_;
  assign new_n4973_ = new_n4321_ & new_n4319_;
  assign new_n4974_ = new_n4320_ | new_n4318_;
  assign new_n4975_ = new_n4317_ & new_n4315_;
  assign new_n4976_ = new_n4316_ | new_n4314_;
  assign new_n4977_ = new_n8742_ & new_n8745_;
  assign new_n4978_ = new_n8748_ | new_n8751_;
  assign new_n4979_ = new_n4977_ & new_n8754_;
  assign new_n4980_ = new_n4978_ | new_n8757_;
  assign new_n4981_ = new_n8742_ & new_n8751_;
  assign new_n4982_ = new_n8748_ | new_n8745_;
  assign new_n4983_ = new_n4981_ & new_n8757_;
  assign new_n4984_ = new_n4982_ | new_n8754_;
  assign new_n4985_ = new_n4984_ & new_n4980_;
  assign new_n4986_ = new_n4983_ | new_n4979_;
  assign new_n4987_ = new_n8749_ & new_n8752_;
  assign new_n4988_ = new_n8743_ | new_n8746_;
  assign new_n4989_ = new_n4987_ & new_n8755_;
  assign new_n4990_ = new_n4988_ | new_n8758_;
  assign new_n4991_ = new_n8749_ & new_n8746_;
  assign new_n4992_ = new_n8743_ | new_n8752_;
  assign new_n4993_ = new_n4991_ & new_n8758_;
  assign new_n4994_ = new_n4992_ | new_n8755_;
  assign new_n4995_ = new_n4994_ & new_n4990_;
  assign new_n4996_ = new_n4993_ | new_n4989_;
  assign new_n4997_ = new_n4995_ & new_n4985_;
  assign new_n4998_ = new_n4996_ | new_n4986_;
  assign new_n4999_ = new_n4997_ & new_n4972_;
  assign new_n5000_ = new_n4998_ & new_n4971_;
  assign new_n5001_ = new_n5000_ | new_n4999_;
  assign new_n5002_ = new_n4372_ & new_n4179_;
  assign new_n5003_ = new_n4373_ | new_n4178_;
  assign new_n5004_ = new_n4374_ & new_n4177_;
  assign new_n5005_ = new_n4375_ | new_n4176_;
  assign new_n5006_ = new_n5005_ & new_n5003_;
  assign new_n5007_ = new_n5004_ | new_n5002_;
  assign new_n5008_ = new_n4403_ & new_n4175_;
  assign new_n5009_ = new_n4402_ | new_n4174_;
  assign new_n5010_ = new_n4370_ & new_n4208_;
  assign new_n5011_ = new_n4371_ | new_n4209_;
  assign new_n5012_ = new_n5011_ & new_n5009_;
  assign new_n5013_ = new_n5010_ | new_n5008_;
  assign new_n5014_ = new_n8759_ & new_n8760_;
  assign new_n5015_ = new_n8761_ | new_n8762_;
  assign new_n5016_ = new_n8761_ & new_n8762_;
  assign new_n5017_ = new_n8759_ | new_n8760_;
  assign new_n5018_ = new_n5017_ & new_n5015_;
  assign new_n5019_ = new_n5016_ | new_n5014_;
  assign new_n5020_ = new_n4313_ & new_n4311_;
  assign new_n5021_ = new_n4312_ | new_n4310_;
  assign new_n5022_ = new_n4309_ & new_n4307_;
  assign new_n5023_ = new_n4308_ | new_n4306_;
  assign new_n5024_ = new_n8764_ & new_n8767_;
  assign new_n5025_ = new_n8770_ | new_n8773_;
  assign new_n5026_ = new_n5024_ & new_n8776_;
  assign new_n5027_ = new_n5025_ | new_n8779_;
  assign new_n5028_ = new_n8764_ & new_n8773_;
  assign new_n5029_ = new_n8770_ | new_n8767_;
  assign new_n5030_ = new_n5028_ & new_n8779_;
  assign new_n5031_ = new_n5029_ | new_n8776_;
  assign new_n5032_ = new_n5031_ & new_n5027_;
  assign new_n5033_ = new_n5030_ | new_n5026_;
  assign new_n5034_ = new_n8771_ & new_n8774_;
  assign new_n5035_ = new_n8765_ | new_n8768_;
  assign new_n5036_ = new_n5034_ & new_n8777_;
  assign new_n5037_ = new_n5035_ | new_n8780_;
  assign new_n5038_ = new_n8771_ & new_n8768_;
  assign new_n5039_ = new_n8765_ | new_n8774_;
  assign new_n5040_ = new_n5038_ & new_n8780_;
  assign new_n5041_ = new_n5039_ | new_n8777_;
  assign new_n5042_ = new_n5041_ & new_n5037_;
  assign new_n5043_ = new_n5040_ | new_n5036_;
  assign new_n5044_ = new_n5042_ & new_n5032_;
  assign new_n5045_ = new_n5043_ | new_n5033_;
  assign new_n5046_ = new_n5044_ & new_n5019_;
  assign new_n5047_ = new_n5045_ & new_n5018_;
  assign new_n5048_ = new_n5047_ | new_n5046_;
  assign new_n5049_ = new_n3853_ | new_n8782_;
  assign new_n5050_ = new_n8602_ | new_n3845_;
  assign new_n5051_ = new_n8603_ | new_n8600_;
  assign new_n5052_ = new_n5051_ | new_n3833_;
  assign new_n5053_ = new_n8603_ | new_n8598_;
  assign new_n5054_ = new_n5053_ | new_n3825_;
  assign new_n5055_ = new_n5054_ | new_n8599_;
  assign new_n5056_ = new_n5050_ & new_n8783_;
  assign new_n5057_ = new_n5056_ & new_n5052_;
  assign new_n5058_ = new_n5057_ & new_n5055_;
  assign new_n5059_ = new_n8604_ | new_n4001_;
  assign new_n5060_ = new_n5059_ & new_n5058_;
  assign new_n5061_ = new_n8613_ | new_n8784_;
  assign new_n5062_ = new_n8614_ | new_n8607_;
  assign new_n5063_ = new_n5062_ | new_n8785_;
  assign new_n5064_ = new_n8614_ | new_n8610_;
  assign new_n5065_ = new_n5064_ | new_n8786_;
  assign new_n5066_ = new_n5065_ | new_n8608_;
  assign new_n5067_ = new_n5061_ & new_n8788_;
  assign new_n5068_ = new_n5067_ & new_n5063_;
  assign new_n5069_ = new_n5068_ & new_n5066_;
  assign new_n5070_ = new_n3850_ & new_n8559_;
  assign new_n5071_ = new_n3851_ | new_n8555_;
  assign new_n5072_ = new_n8648_ & new_n8790_;
  assign new_n5073_ = new_n8653_ | new_n8791_;
  assign new_n5074_ = new_n8619_ & new_n8649_;
  assign new_n5075_ = new_n8629_ | new_n8654_;
  assign new_n5076_ = new_n5074_ & new_n8793_;
  assign new_n5077_ = new_n5075_ | new_n8795_;
  assign new_n5078_ = new_n8638_ & new_n8649_;
  assign new_n5079_ = new_n8643_ | new_n8654_;
  assign new_n5080_ = new_n5078_ & new_n8797_;
  assign new_n5081_ = new_n5079_ | new_n8799_;
  assign new_n5082_ = new_n5080_ & new_n8618_;
  assign new_n5083_ = new_n5081_ | new_n8628_;
  assign new_n5084_ = new_n8658_ & new_n8639_;
  assign new_n5085_ = new_n8663_ | new_n8644_;
  assign new_n5086_ = new_n8800_ & new_n8650_;
  assign new_n5087_ = new_n8801_ | new_n8655_;
  assign new_n5088_ = new_n5086_ & new_n8803_;
  assign new_n5089_ = new_n5087_ | new_n8806_;
  assign new_n5090_ = new_n5088_ & new_n8620_;
  assign new_n5091_ = new_n5089_ | new_n8630_;
  assign new_n5092_ = new_n5073_ & new_n5071_;
  assign new_n5093_ = new_n5072_ | new_n5070_;
  assign new_n5094_ = new_n5092_ & new_n5077_;
  assign new_n5095_ = new_n5093_ | new_n5076_;
  assign new_n5096_ = new_n5094_ & new_n5083_;
  assign new_n5097_ = new_n5095_ | new_n5082_;
  assign new_n5098_ = new_n5096_ & new_n5091_;
  assign new_n5099_ = new_n5097_ | new_n5090_;
  assign new_n5100_ = new_n8808_ | new_n8667_;
  assign new_n5101_ = new_n5100_ & new_n5069_;
  assign new_n5102_ = new_n8683_ | new_n8809_;
  assign new_n5103_ = new_n8682_ | new_n8677_;
  assign new_n5104_ = new_n5103_ | new_n8810_;
  assign new_n5105_ = new_n8684_ | new_n8680_;
  assign new_n5106_ = new_n5105_ | new_n8811_;
  assign new_n5107_ = new_n5106_ | new_n8678_;
  assign new_n5108_ = new_n5102_ & new_n8783_;
  assign new_n5109_ = new_n5108_ & new_n5104_;
  assign new_n5110_ = new_n5109_ & new_n5107_;
  assign new_n5111_ = new_n3848_ & new_n8568_;
  assign new_n5112_ = new_n3849_ | new_n8564_;
  assign new_n5113_ = new_n8717_ & new_n8812_;
  assign new_n5114_ = new_n8722_ | new_n8813_;
  assign new_n5115_ = new_n8718_ & new_n8688_;
  assign new_n5116_ = new_n8723_ | new_n8698_;
  assign new_n5117_ = new_n5115_ & new_n8815_;
  assign new_n5118_ = new_n5116_ | new_n8817_;
  assign new_n5119_ = new_n8718_ & new_n8707_;
  assign new_n5120_ = new_n8723_ | new_n8712_;
  assign new_n5121_ = new_n5119_ & new_n8819_;
  assign new_n5122_ = new_n5120_ | new_n8821_;
  assign new_n5123_ = new_n5121_ & new_n8687_;
  assign new_n5124_ = new_n5122_ | new_n8697_;
  assign new_n5125_ = new_n8727_ & new_n8708_;
  assign new_n5126_ = new_n8732_ | new_n8713_;
  assign new_n5127_ = new_n8822_ & new_n8719_;
  assign new_n5128_ = new_n8823_ | new_n8724_;
  assign new_n5129_ = new_n5127_ & new_n8825_;
  assign new_n5130_ = new_n5128_ | new_n8828_;
  assign new_n5131_ = new_n5129_ & new_n8689_;
  assign new_n5132_ = new_n5130_ | new_n8699_;
  assign new_n5133_ = new_n5114_ & new_n5112_;
  assign new_n5134_ = new_n5113_ | new_n5111_;
  assign new_n5135_ = new_n5133_ & new_n5118_;
  assign new_n5136_ = new_n5134_ | new_n5117_;
  assign new_n5137_ = new_n5135_ & new_n5124_;
  assign new_n5138_ = new_n5136_ | new_n5123_;
  assign new_n5139_ = new_n5137_ & new_n5132_;
  assign new_n5140_ = new_n5138_ | new_n5131_;
  assign new_n5141_ = new_n8830_ | new_n8736_;
  assign new_n5142_ = new_n5141_ & new_n5110_;
  assign new_n5143_ = new_n8672_ | new_n3846_;
  assign new_n5144_ = new_n8673_ | new_n8670_;
  assign new_n5145_ = new_n5144_ | new_n3835_;
  assign new_n5146_ = new_n8673_ | new_n8668_;
  assign new_n5147_ = new_n5146_ | new_n3827_;
  assign new_n5148_ = new_n5147_ | new_n8669_;
  assign new_n5149_ = new_n5143_ & new_n8788_;
  assign new_n5150_ = new_n5149_ & new_n5145_;
  assign new_n5151_ = new_n5150_ & new_n5148_;
  assign new_n5152_ = new_n8674_ | new_n4003_;
  assign new_n5153_ = new_n5152_ & new_n5151_;
  assign new_n5154_ = new_n8831_ | new_n3516_;
  assign new_n5155_ = new_n8832_ | new_n3517_;
  assign new_n5156_ = new_n5155_ & new_n5154_;
  assign new_n5157_ = new_n5156_ & new_n8838_;
  assign new_n5158_ = new_n5157_ & new_n8878_;
  assign new_n5159_ = new_n8635_ & new_n8914_;
  assign new_n5160_ = new_n8625_ & new_n8916_;
  assign new_n5161_ = new_n5160_ | new_n5159_;
  assign new_n5162_ = new_n8917_ & new_n8922_;
  assign new_n5163_ = new_n5162_ & new_n8878_;
  assign new_n5164_ = new_n8838_ & new_n3162_;
  assign new_n5165_ = new_n5164_ & new_n8945_;
  assign new_n5166_ = new_n5163_ | new_n5158_;
  assign new_n5167_ = new_n5166_ | new_n5165_;
  assign new_n5168_ = new_n8561_ & new_n8839_;
  assign new_n5169_ = new_n5168_ & new_n8879_;
  assign new_n5170_ = new_n8624_ & new_n8914_;
  assign new_n5171_ = new_n8634_ | new_n8916_;
  assign new_n5172_ = new_n8965_ & new_n8806_;
  assign new_n5173_ = new_n8967_ | new_n8803_;
  assign new_n5174_ = new_n5172_ & new_n8664_;
  assign new_n5175_ = new_n5173_ & new_n8659_;
  assign new_n5176_ = new_n5175_ | new_n5174_;
  assign new_n5177_ = new_n8968_ & new_n8922_;
  assign new_n5178_ = new_n5177_ & new_n8879_;
  assign new_n5179_ = new_n8839_ & new_n3146_;
  assign new_n5180_ = new_n5179_ & new_n8945_;
  assign new_n5181_ = new_n5178_ | new_n5169_;
  assign new_n5182_ = new_n5181_ | new_n5180_;
  assign new_n5183_ = new_n8595_ & new_n8841_;
  assign new_n5184_ = new_n5183_ & new_n8881_;
  assign new_n5185_ = new_n8704_ & new_n8970_;
  assign new_n5186_ = new_n8694_ & new_n8972_;
  assign new_n5187_ = new_n5186_ | new_n5185_;
  assign new_n5188_ = new_n8973_ & new_n8923_;
  assign new_n5189_ = new_n5188_ & new_n8881_;
  assign new_n5190_ = new_n8841_ & new_n3066_;
  assign new_n5191_ = new_n5190_ & new_n8946_;
  assign new_n5192_ = new_n5189_ | new_n5184_;
  assign new_n5193_ = new_n5192_ | new_n5191_;
  assign new_n5194_ = new_n8974_ & new_n8975_;
  assign new_n5195_ = new_n8976_ | new_n8977_;
  assign new_n5196_ = new_n8976_ & new_n8977_;
  assign new_n5197_ = new_n8974_ | new_n8975_;
  assign new_n5198_ = new_n5197_ & new_n5195_;
  assign new_n5199_ = new_n5196_ | new_n5194_;
  assign new_n5200_ = new_n4936_ & new_n8913_;
  assign new_n5201_ = new_n8666_ | new_n8915_;
  assign new_n5202_ = new_n5201_ & new_n8808_;
  assign new_n5203_ = new_n5200_ | new_n5099_;
  assign new_n5204_ = new_n8980_ & new_n5198_;
  assign new_n5205_ = new_n8984_ | new_n5199_;
  assign new_n5206_ = new_n4331_ & new_n8784_;
  assign new_n5207_ = new_n4330_ | new_n4205_;
  assign new_n5208_ = new_n5206_ & new_n4335_;
  assign new_n5209_ = new_n5207_ | new_n4334_;
  assign new_n5210_ = new_n5208_ & new_n4353_;
  assign new_n5211_ = new_n5209_ | new_n4352_;
  assign new_n5212_ = new_n8986_ & new_n8615_;
  assign new_n5213_ = new_n8987_ | new_n8988_;
  assign new_n5214_ = new_n8987_ & new_n8988_;
  assign new_n5215_ = new_n8986_ | new_n8615_;
  assign new_n5216_ = new_n5215_ & new_n5213_;
  assign new_n5217_ = new_n5214_ | new_n5212_;
  assign new_n5218_ = new_n5217_ & new_n8984_;
  assign new_n5219_ = new_n5216_ | new_n8980_;
  assign new_n5220_ = new_n5219_ & new_n5205_;
  assign new_n5221_ = new_n5218_ | new_n5204_;
  assign new_n5222_ = new_n8991_ & new_n8997_;
  assign new_n5223_ = new_n5222_ & new_n9016_;
  assign new_n5224_ = new_n9033_ & new_n9039_;
  assign new_n5225_ = new_n5224_ & new_n9016_;
  assign new_n5226_ = new_n8997_ & new_n9054_;
  assign new_n5227_ = new_n5226_ & new_n9059_;
  assign new_n5228_ = new_n9039_ & new_n9074_;
  assign new_n5229_ = new_n5228_ & new_n9059_;
  assign new_n5230_ = new_n5225_ | new_n5223_;
  assign new_n5231_ = new_n5230_ | new_n5227_;
  assign new_n5232_ = new_n5231_ | new_n5229_;
  assign new_n5233_ = new_n8563_ & new_n8842_;
  assign new_n5234_ = new_n5233_ & new_n8882_;
  assign new_n5235_ = new_n8620_ & new_n8793_;
  assign new_n5236_ = new_n8630_ | new_n8795_;
  assign new_n5237_ = new_n8639_ & new_n8797_;
  assign new_n5238_ = new_n8644_ | new_n8799_;
  assign new_n5239_ = new_n9075_ & new_n8622_;
  assign new_n5240_ = new_n9076_ | new_n8632_;
  assign new_n5241_ = new_n8800_ & new_n8804_;
  assign new_n5242_ = new_n8801_ | new_n8807_;
  assign new_n5243_ = new_n9077_ & new_n8622_;
  assign new_n5244_ = new_n9078_ | new_n8632_;
  assign new_n5245_ = new_n8967_ & new_n8640_;
  assign new_n5246_ = new_n8965_ | new_n8645_;
  assign new_n5247_ = new_n5245_ & new_n8659_;
  assign new_n5248_ = new_n5246_ | new_n8664_;
  assign new_n5249_ = new_n9079_ & new_n8623_;
  assign new_n5250_ = new_n9080_ | new_n8633_;
  assign new_n5251_ = new_n5236_ & new_n8791_;
  assign new_n5252_ = new_n5235_ | new_n8790_;
  assign new_n5253_ = new_n5251_ & new_n5240_;
  assign new_n5254_ = new_n5252_ | new_n5239_;
  assign new_n5255_ = new_n5253_ & new_n5244_;
  assign new_n5256_ = new_n5254_ | new_n5243_;
  assign new_n5257_ = new_n5255_ & new_n5250_;
  assign new_n5258_ = new_n5256_ | new_n5249_;
  assign new_n5259_ = new_n5257_ & new_n8655_;
  assign new_n5260_ = new_n5258_ & new_n8650_;
  assign new_n5261_ = new_n5260_ | new_n5259_;
  assign new_n5262_ = new_n9081_ & new_n8923_;
  assign new_n5263_ = new_n5262_ & new_n8882_;
  assign new_n5264_ = new_n8842_ & new_n2834_;
  assign new_n5265_ = new_n5264_ & new_n8946_;
  assign new_n5266_ = new_n5263_ | new_n5234_;
  assign new_n5267_ = new_n5266_ | new_n5265_;
  assign new_n5268_ = new_n8562_ & new_n8845_;
  assign new_n5269_ = new_n5268_ & new_n8885_;
  assign new_n5270_ = new_n9076_ & new_n8794_;
  assign new_n5271_ = new_n9075_ | new_n8792_;
  assign new_n5272_ = new_n5270_ & new_n9078_;
  assign new_n5273_ = new_n5271_ | new_n9077_;
  assign new_n5274_ = new_n5272_ & new_n9080_;
  assign new_n5275_ = new_n5273_ | new_n9079_;
  assign new_n5276_ = new_n5274_ & new_n8633_;
  assign new_n5277_ = new_n5275_ & new_n8623_;
  assign new_n5278_ = new_n5277_ | new_n5276_;
  assign new_n5279_ = new_n9082_ & new_n8925_;
  assign new_n5280_ = new_n5279_ & new_n8885_;
  assign new_n5281_ = new_n8845_ & new_n3154_;
  assign new_n5282_ = new_n5281_ & new_n8948_;
  assign new_n5283_ = new_n5280_ | new_n5269_;
  assign new_n5284_ = new_n5283_ | new_n5282_;
  assign new_n5285_ = new_n8560_ & new_n8846_;
  assign new_n5286_ = new_n5285_ & new_n8886_;
  assign new_n5287_ = new_n8660_ & new_n8804_;
  assign new_n5288_ = new_n8665_ | new_n8807_;
  assign new_n5289_ = new_n8966_ & new_n8660_;
  assign new_n5290_ = new_n8964_ | new_n8665_;
  assign new_n5291_ = new_n5288_ & new_n8798_;
  assign new_n5292_ = new_n5287_ | new_n8796_;
  assign new_n5293_ = new_n5291_ & new_n5290_;
  assign new_n5294_ = new_n5292_ | new_n5289_;
  assign new_n5295_ = new_n5293_ & new_n8645_;
  assign new_n5296_ = new_n5294_ & new_n8640_;
  assign new_n5297_ = new_n5296_ | new_n5295_;
  assign new_n5298_ = new_n9083_ & new_n8925_;
  assign new_n5299_ = new_n5298_ & new_n8886_;
  assign new_n5300_ = new_n8846_ & new_n3082_;
  assign new_n5301_ = new_n5300_ & new_n8948_;
  assign new_n5302_ = new_n5299_ | new_n5286_;
  assign new_n5303_ = new_n5302_ | new_n5301_;
  assign new_n5304_ = new_n8991_ & new_n9088_;
  assign new_n5305_ = new_n5304_ & new_n9107_;
  assign new_n5306_ = new_n9033_ & new_n9126_;
  assign new_n5307_ = new_n5306_ & new_n9107_;
  assign new_n5308_ = new_n9088_ & new_n9054_;
  assign new_n5309_ = new_n5308_ & new_n9145_;
  assign new_n5310_ = new_n9126_ & new_n9074_;
  assign new_n5311_ = new_n5310_ & new_n9145_;
  assign new_n5312_ = new_n5307_ | new_n5305_;
  assign new_n5313_ = new_n5312_ | new_n5309_;
  assign new_n5314_ = new_n5313_ | new_n5311_;
  assign new_n5315_ = new_n8579_ & new_n8848_;
  assign new_n5316_ = new_n5315_ & new_n8888_;
  assign new_n5317_ = new_n8689_ & new_n8815_;
  assign new_n5318_ = new_n8699_ | new_n8817_;
  assign new_n5319_ = new_n8708_ & new_n8819_;
  assign new_n5320_ = new_n8713_ | new_n8821_;
  assign new_n5321_ = new_n9160_ & new_n8691_;
  assign new_n5322_ = new_n9161_ | new_n8701_;
  assign new_n5323_ = new_n8822_ & new_n8825_;
  assign new_n5324_ = new_n8823_ | new_n8828_;
  assign new_n5325_ = new_n9162_ & new_n8691_;
  assign new_n5326_ = new_n9163_ | new_n8701_;
  assign new_n5327_ = new_n8693_ & new_n8970_;
  assign new_n5328_ = new_n8703_ | new_n8972_;
  assign new_n5329_ = new_n9165_ & new_n8709_;
  assign new_n5330_ = new_n9167_ | new_n8714_;
  assign new_n5331_ = new_n5329_ & new_n8728_;
  assign new_n5332_ = new_n5330_ | new_n8733_;
  assign new_n5333_ = new_n9168_ & new_n8692_;
  assign new_n5334_ = new_n9169_ | new_n8702_;
  assign new_n5335_ = new_n5318_ & new_n8813_;
  assign new_n5336_ = new_n5317_ | new_n8812_;
  assign new_n5337_ = new_n5335_ & new_n5322_;
  assign new_n5338_ = new_n5336_ | new_n5321_;
  assign new_n5339_ = new_n5337_ & new_n5326_;
  assign new_n5340_ = new_n5338_ | new_n5325_;
  assign new_n5341_ = new_n5339_ & new_n5334_;
  assign new_n5342_ = new_n5340_ | new_n5333_;
  assign new_n5343_ = new_n5341_ & new_n8724_;
  assign new_n5344_ = new_n5342_ & new_n8719_;
  assign new_n5345_ = new_n5344_ | new_n5343_;
  assign new_n5346_ = new_n9170_ & new_n8926_;
  assign new_n5347_ = new_n5346_ & new_n8888_;
  assign new_n5348_ = new_n8848_ & new_n3106_;
  assign new_n5349_ = new_n5348_ & new_n8949_;
  assign new_n5350_ = new_n5347_ | new_n5316_;
  assign new_n5351_ = new_n5350_ | new_n5349_;
  assign new_n5352_ = new_n8597_ & new_n8849_;
  assign new_n5353_ = new_n5352_ & new_n8889_;
  assign new_n5354_ = new_n9161_ & new_n8816_;
  assign new_n5355_ = new_n9160_ | new_n8814_;
  assign new_n5356_ = new_n5354_ & new_n9163_;
  assign new_n5357_ = new_n5355_ | new_n9162_;
  assign new_n5358_ = new_n5356_ & new_n9169_;
  assign new_n5359_ = new_n5357_ | new_n9168_;
  assign new_n5360_ = new_n5358_ & new_n8702_;
  assign new_n5361_ = new_n5359_ & new_n8692_;
  assign new_n5362_ = new_n5361_ | new_n5360_;
  assign new_n5363_ = new_n9171_ & new_n8926_;
  assign new_n5364_ = new_n5363_ & new_n8889_;
  assign new_n5365_ = new_n8849_ & new_n3138_;
  assign new_n5366_ = new_n5365_ & new_n8949_;
  assign new_n5367_ = new_n5364_ | new_n5353_;
  assign new_n5368_ = new_n5367_ | new_n5366_;
  assign new_n5369_ = new_n8596_ & new_n8853_;
  assign new_n5370_ = new_n5369_ & new_n8893_;
  assign new_n5371_ = new_n8728_ & new_n8826_;
  assign new_n5372_ = new_n8733_ | new_n8829_;
  assign new_n5373_ = new_n9165_ & new_n8729_;
  assign new_n5374_ = new_n9167_ | new_n8734_;
  assign new_n5375_ = new_n5372_ & new_n8820_;
  assign new_n5376_ = new_n5371_ | new_n8818_;
  assign new_n5377_ = new_n5375_ & new_n5374_;
  assign new_n5378_ = new_n5376_ | new_n5373_;
  assign new_n5379_ = new_n5377_ & new_n8714_;
  assign new_n5380_ = new_n5378_ & new_n8709_;
  assign new_n5381_ = new_n5380_ | new_n5379_;
  assign new_n5382_ = new_n9172_ & new_n8929_;
  assign new_n5383_ = new_n5382_ & new_n8893_;
  assign new_n5384_ = new_n8853_ & new_n3130_;
  assign new_n5385_ = new_n5384_ & new_n8952_;
  assign new_n5386_ = new_n5383_ | new_n5370_;
  assign new_n5387_ = new_n5386_ | new_n5385_;
  assign new_n5388_ = new_n8594_ & new_n8852_;
  assign new_n5389_ = new_n5388_ & new_n8892_;
  assign new_n5390_ = new_n9166_ & new_n8829_;
  assign new_n5391_ = new_n9164_ | new_n8826_;
  assign new_n5392_ = new_n5390_ & new_n8734_;
  assign new_n5393_ = new_n5391_ & new_n8729_;
  assign new_n5394_ = new_n5393_ | new_n5392_;
  assign new_n5395_ = new_n9173_ & new_n8929_;
  assign new_n5396_ = new_n5395_ & new_n8894_;
  assign new_n5397_ = new_n8854_ & new_n3122_;
  assign new_n5398_ = new_n5397_ & new_n8952_;
  assign new_n5399_ = new_n5396_ | new_n5389_;
  assign new_n5400_ = new_n5399_ | new_n5398_;
  assign new_n5401_ = new_n4394_ & new_n4203_;
  assign new_n5402_ = new_n4395_ | new_n4202_;
  assign new_n5403_ = new_n4396_ & new_n4201_;
  assign new_n5404_ = new_n4397_ | new_n4200_;
  assign new_n5405_ = new_n5404_ & new_n5402_;
  assign new_n5406_ = new_n5403_ | new_n5401_;
  assign new_n5407_ = new_n4406_ & new_n4207_;
  assign new_n5408_ = new_n4407_ | new_n4206_;
  assign new_n5409_ = new_n4400_ & new_n4213_;
  assign new_n5410_ = new_n4401_ | new_n4212_;
  assign new_n5411_ = new_n5410_ & new_n5408_;
  assign new_n5412_ = new_n5409_ | new_n5407_;
  assign new_n5413_ = new_n9174_ & new_n9175_;
  assign new_n5414_ = new_n9176_ | new_n9177_;
  assign new_n5415_ = new_n9176_ & new_n9177_;
  assign new_n5416_ = new_n9174_ | new_n9175_;
  assign new_n5417_ = new_n5416_ & new_n5414_;
  assign new_n5418_ = new_n5415_ | new_n5413_;
  assign new_n5419_ = new_n4341_ & new_n4339_;
  assign new_n5420_ = new_n4340_ | new_n4338_;
  assign new_n5421_ = new_n4357_ & new_n4342_;
  assign new_n5422_ = new_n4356_ | new_n4343_;
  assign new_n5423_ = new_n9179_ & new_n9182_;
  assign new_n5424_ = new_n9185_ | new_n9188_;
  assign new_n5425_ = new_n5423_ & new_n9191_;
  assign new_n5426_ = new_n5424_ | new_n9194_;
  assign new_n5427_ = new_n9179_ & new_n9188_;
  assign new_n5428_ = new_n9185_ | new_n9182_;
  assign new_n5429_ = new_n5427_ & new_n9194_;
  assign new_n5430_ = new_n5428_ | new_n9191_;
  assign new_n5431_ = new_n5430_ & new_n5426_;
  assign new_n5432_ = new_n5429_ | new_n5425_;
  assign new_n5433_ = new_n9186_ & new_n9189_;
  assign new_n5434_ = new_n9180_ | new_n9183_;
  assign new_n5435_ = new_n5433_ & new_n9192_;
  assign new_n5436_ = new_n5434_ | new_n9195_;
  assign new_n5437_ = new_n9186_ & new_n9183_;
  assign new_n5438_ = new_n9180_ | new_n9189_;
  assign new_n5439_ = new_n5437_ & new_n9195_;
  assign new_n5440_ = new_n5438_ | new_n9192_;
  assign new_n5441_ = new_n5440_ & new_n5436_;
  assign new_n5442_ = new_n5439_ | new_n5435_;
  assign new_n5443_ = new_n5441_ & new_n5431_;
  assign new_n5444_ = new_n5442_ | new_n5432_;
  assign new_n5445_ = new_n5443_ & new_n5418_;
  assign new_n5446_ = new_n5444_ & new_n5417_;
  assign new_n5447_ = new_n5446_ | new_n5445_;
  assign new_n5448_ = new_n4388_ & new_n4197_;
  assign new_n5449_ = new_n4389_ | new_n4196_;
  assign new_n5450_ = new_n4390_ & new_n4195_;
  assign new_n5451_ = new_n4391_ | new_n4194_;
  assign new_n5452_ = new_n5451_ & new_n5449_;
  assign new_n5453_ = new_n5450_ | new_n5448_;
  assign new_n5454_ = new_n4392_ & new_n4193_;
  assign new_n5455_ = new_n4393_ | new_n4192_;
  assign new_n5456_ = new_n4386_ & new_n4199_;
  assign new_n5457_ = new_n4387_ | new_n4198_;
  assign new_n5458_ = new_n5457_ & new_n5455_;
  assign new_n5459_ = new_n5456_ | new_n5454_;
  assign new_n5460_ = new_n9196_ & new_n9197_;
  assign new_n5461_ = new_n9198_ | new_n9199_;
  assign new_n5462_ = new_n9198_ & new_n9199_;
  assign new_n5463_ = new_n9196_ | new_n9197_;
  assign new_n5464_ = new_n5463_ & new_n5461_;
  assign new_n5465_ = new_n5462_ | new_n5460_;
  assign new_n5466_ = new_n4355_ & new_n4347_;
  assign new_n5467_ = new_n4354_ | new_n4346_;
  assign new_n5468_ = new_n4349_ & new_n4345_;
  assign new_n5469_ = new_n4348_ | new_n4344_;
  assign new_n5470_ = new_n9201_ & new_n9204_;
  assign new_n5471_ = new_n9207_ | new_n9210_;
  assign new_n5472_ = new_n5470_ & new_n9213_;
  assign new_n5473_ = new_n5471_ | new_n9216_;
  assign new_n5474_ = new_n9201_ & new_n9210_;
  assign new_n5475_ = new_n9207_ | new_n9204_;
  assign new_n5476_ = new_n5474_ & new_n9216_;
  assign new_n5477_ = new_n5475_ | new_n9213_;
  assign new_n5478_ = new_n5477_ & new_n5473_;
  assign new_n5479_ = new_n5476_ | new_n5472_;
  assign new_n5480_ = new_n9208_ & new_n9211_;
  assign new_n5481_ = new_n9202_ | new_n9205_;
  assign new_n5482_ = new_n5480_ & new_n9214_;
  assign new_n5483_ = new_n5481_ | new_n9217_;
  assign new_n5484_ = new_n9208_ & new_n9205_;
  assign new_n5485_ = new_n9202_ | new_n9211_;
  assign new_n5486_ = new_n5484_ & new_n9217_;
  assign new_n5487_ = new_n5485_ | new_n9214_;
  assign new_n5488_ = new_n5487_ & new_n5483_;
  assign new_n5489_ = new_n5486_ | new_n5482_;
  assign new_n5490_ = new_n5488_ & new_n5478_;
  assign new_n5491_ = new_n5489_ | new_n5479_;
  assign new_n5492_ = new_n5490_ & new_n5465_;
  assign new_n5493_ = new_n5491_ & new_n5464_;
  assign new_n5494_ = new_n5493_ | new_n5492_;
  assign new_n5495_ = new_n4952_ & new_n8969_;
  assign new_n5496_ = new_n8735_ | new_n8971_;
  assign new_n5497_ = new_n5496_ & new_n8830_;
  assign new_n5498_ = new_n5495_ | new_n5140_;
  assign new_n5499_ = new_n9219_ & new_n4222_;
  assign new_n5500_ = new_n9222_ & new_n8675_;
  assign new_n5501_ = new_n5500_ | new_n5499_;
  assign new_n5502_ = new_n8679_ & new_n4104_;
  assign new_n5503_ = new_n4120_ & new_n8811_;
  assign new_n5504_ = new_n5503_ | new_n5502_;
  assign new_n5505_ = new_n5504_ & new_n9219_;
  assign new_n5506_ = new_n4364_ | new_n4271_;
  assign new_n5507_ = new_n4365_ | new_n4270_;
  assign new_n5508_ = new_n5507_ & new_n5506_;
  assign new_n5509_ = new_n5508_ & new_n9222_;
  assign new_n5510_ = new_n5509_ | new_n5505_;
  assign new_n5511_ = new_n4360_ | new_n4329_;
  assign new_n5512_ = new_n4361_ | new_n4328_;
  assign new_n5513_ = new_n5512_ & new_n5511_;
  assign new_n5514_ = new_n5513_ & new_n9220_;
  assign new_n5515_ = new_n4325_ & new_n8810_;
  assign new_n5516_ = new_n4324_ | new_n4106_;
  assign new_n5517_ = new_n5515_ & new_n4363_;
  assign new_n5518_ = new_n5516_ | new_n4362_;
  assign new_n5519_ = new_n5517_ & new_n8678_;
  assign new_n5520_ = new_n5518_ & new_n4118_;
  assign new_n5521_ = new_n5520_ | new_n5519_;
  assign new_n5522_ = new_n5521_ & new_n9223_;
  assign new_n5523_ = new_n5522_ | new_n5514_;
  assign new_n5524_ = new_n4444_ | new_n4385_;
  assign new_n5525_ = new_n4445_ | new_n4384_;
  assign new_n5526_ = new_n5525_ & new_n5524_;
  assign new_n5527_ = new_n5526_ & new_n9220_;
  assign new_n5528_ = new_n4327_ & new_n8809_;
  assign new_n5529_ = new_n4326_ | new_n4190_;
  assign new_n5530_ = new_n5528_ & new_n4323_;
  assign new_n5531_ = new_n5529_ | new_n4322_;
  assign new_n5532_ = new_n5530_ & new_n4359_;
  assign new_n5533_ = new_n5531_ | new_n4358_;
  assign new_n5534_ = new_n5532_ & new_n8684_;
  assign new_n5535_ = new_n5533_ & new_n4224_;
  assign new_n5536_ = new_n5535_ | new_n5534_;
  assign new_n5537_ = new_n5536_ & new_n9223_;
  assign new_n5538_ = new_n5537_ | new_n5527_;
  assign new_n5539_ = new_n9173_ | new_n8973_;
  assign new_n5540_ = new_n5539_ | new_n9172_;
  assign new_n5541_ = new_n5540_ | new_n9171_;
  assign new_n5542_ = new_n5541_ | new_n9170_;
  assign new_n5543_ = new_n5542_ | new_n9224_;
  assign new_n5544_ = new_n5543_ | new_n9225_;
  assign new_n5545_ = new_n5544_ | new_n9226_;
  assign new_n5546_ = new_n5545_ | new_n9227_;
  assign new_n5547_ = new_n8979_ & new_n4226_;
  assign new_n5548_ = new_n8983_ & new_n8605_;
  assign new_n5549_ = new_n5548_ | new_n5547_;
  assign new_n5550_ = new_n8609_ & new_n4110_;
  assign new_n5551_ = new_n4122_ & new_n8786_;
  assign new_n5552_ = new_n5551_ | new_n5550_;
  assign new_n5553_ = new_n5552_ & new_n8981_;
  assign new_n5554_ = new_n4368_ | new_n4273_;
  assign new_n5555_ = new_n4369_ | new_n4272_;
  assign new_n5556_ = new_n5555_ & new_n5554_;
  assign new_n5557_ = new_n5556_ & new_n8985_;
  assign new_n5558_ = new_n5557_ | new_n5553_;
  assign new_n5559_ = new_n4351_ | new_n4333_;
  assign new_n5560_ = new_n4350_ | new_n4332_;
  assign new_n5561_ = new_n5560_ & new_n5559_;
  assign new_n5562_ = new_n5561_ & new_n8981_;
  assign new_n5563_ = new_n4337_ & new_n8785_;
  assign new_n5564_ = new_n4336_ | new_n4108_;
  assign new_n5565_ = new_n5563_ & new_n4367_;
  assign new_n5566_ = new_n5564_ | new_n4366_;
  assign new_n5567_ = new_n5565_ & new_n8608_;
  assign new_n5568_ = new_n5566_ & new_n4113_;
  assign new_n5569_ = new_n5568_ | new_n5567_;
  assign new_n5570_ = new_n5569_ & new_n8985_;
  assign new_n5571_ = new_n5570_ | new_n5562_;
  assign new_n5572_ = new_n8968_ | new_n8917_;
  assign new_n5573_ = new_n5572_ | new_n9083_;
  assign new_n5574_ = new_n5573_ | new_n9082_;
  assign new_n5575_ = new_n5574_ | new_n9081_;
  assign new_n5576_ = new_n5575_ | new_n9228_;
  assign new_n5577_ = new_n5576_ | new_n9229_;
  assign new_n5578_ = new_n5577_ | new_n9230_;
  assign new_n5579_ = new_n5578_ | new_n9232_;
  assign new_n5580_ = new_n8990_ & new_n9238_;
  assign new_n5581_ = new_n5580_ & new_n9257_;
  assign new_n5582_ = new_n9032_ & new_n9276_;
  assign new_n5583_ = new_n5582_ & new_n9257_;
  assign new_n5584_ = new_n9238_ & new_n9291_;
  assign new_n5585_ = new_n5584_ & new_n9296_;
  assign new_n5586_ = new_n9276_ & new_n9311_;
  assign new_n5587_ = new_n5586_ & new_n9296_;
  assign new_n5588_ = new_n5583_ | new_n5581_;
  assign new_n5589_ = new_n5588_ | new_n5585_;
  assign new_n5590_ = new_n5589_ | new_n5587_;
  assign new_n5591_ = new_n5590_ & new_n9316_;
  assign new_n5592_ = new_n8992_ & new_n9336_;
  assign new_n5593_ = new_n5592_ & new_n9355_;
  assign new_n5594_ = new_n9034_ & new_n9374_;
  assign new_n5595_ = new_n5594_ & new_n9355_;
  assign new_n5596_ = new_n9336_ & new_n9291_;
  assign new_n5597_ = new_n5596_ & new_n9393_;
  assign new_n5598_ = new_n9374_ & new_n9311_;
  assign new_n5599_ = new_n5598_ & new_n9393_;
  assign new_n5600_ = new_n5595_ | new_n5593_;
  assign new_n5601_ = new_n5600_ | new_n5597_;
  assign new_n5602_ = new_n5601_ | new_n5599_;
  assign new_n5603_ = new_n5602_ & new_n9316_;
  assign new_n5604_ = new_n9410_ & new_n8998_;
  assign new_n5605_ = new_n5604_ & new_n9017_;
  assign new_n5606_ = new_n9414_ & new_n9040_;
  assign new_n5607_ = new_n5606_ & new_n9017_;
  assign new_n5608_ = new_n8998_ & new_n9416_;
  assign new_n5609_ = new_n5608_ & new_n9060_;
  assign new_n5610_ = new_n9040_ & new_n9417_;
  assign new_n5611_ = new_n5610_ & new_n9060_;
  assign new_n5612_ = new_n5607_ | new_n5605_;
  assign new_n5613_ = new_n5612_ | new_n5609_;
  assign new_n5614_ = new_n5613_ | new_n5611_;
  assign new_n5615_ = new_n9420_ & new_n9000_;
  assign new_n5616_ = new_n5615_ & new_n9019_;
  assign new_n5617_ = new_n9424_ & new_n9042_;
  assign new_n5618_ = new_n5617_ & new_n9019_;
  assign new_n5619_ = new_n9000_ & new_n9426_;
  assign new_n5620_ = new_n5619_ & new_n9062_;
  assign new_n5621_ = new_n9042_ & new_n9427_;
  assign new_n5622_ = new_n5621_ & new_n9062_;
  assign new_n5623_ = new_n5618_ | new_n5616_;
  assign new_n5624_ = new_n5623_ | new_n5620_;
  assign new_n5625_ = new_n5624_ | new_n5622_;
  assign new_n5626_ = new_n9430_ & new_n9001_;
  assign new_n5627_ = new_n5626_ & new_n9020_;
  assign new_n5628_ = new_n9434_ & new_n9043_;
  assign new_n5629_ = new_n5628_ & new_n9020_;
  assign new_n5630_ = new_n9001_ & new_n9436_;
  assign new_n5631_ = new_n5630_ & new_n9063_;
  assign new_n5632_ = new_n9043_ & new_n9437_;
  assign new_n5633_ = new_n5632_ & new_n9063_;
  assign new_n5634_ = new_n5629_ | new_n5627_;
  assign new_n5635_ = new_n5634_ | new_n5631_;
  assign new_n5636_ = new_n5635_ | new_n5633_;
  assign new_n5637_ = new_n9440_ & new_n9003_;
  assign new_n5638_ = new_n5637_ & new_n9022_;
  assign new_n5639_ = new_n9444_ & new_n9045_;
  assign new_n5640_ = new_n5639_ & new_n9022_;
  assign new_n5641_ = new_n9003_ & new_n9446_;
  assign new_n5642_ = new_n5641_ & new_n9065_;
  assign new_n5643_ = new_n9045_ & new_n9447_;
  assign new_n5644_ = new_n5643_ & new_n9065_;
  assign new_n5645_ = new_n5640_ | new_n5638_;
  assign new_n5646_ = new_n5645_ | new_n5642_;
  assign new_n5647_ = new_n5646_ | new_n5644_;
  assign new_n5648_ = new_n9410_ & new_n9089_;
  assign new_n5649_ = new_n5648_ & new_n9108_;
  assign new_n5650_ = new_n9414_ & new_n9127_;
  assign new_n5651_ = new_n5650_ & new_n9108_;
  assign new_n5652_ = new_n9089_ & new_n9416_;
  assign new_n5653_ = new_n5652_ & new_n9146_;
  assign new_n5654_ = new_n9127_ & new_n9417_;
  assign new_n5655_ = new_n5654_ & new_n9146_;
  assign new_n5656_ = new_n5651_ | new_n5649_;
  assign new_n5657_ = new_n5656_ | new_n5653_;
  assign new_n5658_ = new_n5657_ | new_n5655_;
  assign new_n5659_ = new_n9420_ & new_n9091_;
  assign new_n5660_ = new_n5659_ & new_n9110_;
  assign new_n5661_ = new_n9424_ & new_n9129_;
  assign new_n5662_ = new_n5661_ & new_n9110_;
  assign new_n5663_ = new_n9091_ & new_n9426_;
  assign new_n5664_ = new_n5663_ & new_n9148_;
  assign new_n5665_ = new_n9129_ & new_n9427_;
  assign new_n5666_ = new_n5665_ & new_n9148_;
  assign new_n5667_ = new_n5662_ | new_n5660_;
  assign new_n5668_ = new_n5667_ | new_n5664_;
  assign new_n5669_ = new_n5668_ | new_n5666_;
  assign new_n5670_ = new_n9430_ & new_n9092_;
  assign new_n5671_ = new_n5670_ & new_n9111_;
  assign new_n5672_ = new_n9434_ & new_n9130_;
  assign new_n5673_ = new_n5672_ & new_n9111_;
  assign new_n5674_ = new_n9092_ & new_n9436_;
  assign new_n5675_ = new_n5674_ & new_n9149_;
  assign new_n5676_ = new_n9130_ & new_n9437_;
  assign new_n5677_ = new_n5676_ & new_n9149_;
  assign new_n5678_ = new_n5673_ | new_n5671_;
  assign new_n5679_ = new_n5678_ | new_n5675_;
  assign new_n5680_ = new_n5679_ | new_n5677_;
  assign new_n5681_ = new_n9440_ & new_n9094_;
  assign new_n5682_ = new_n5681_ & new_n9113_;
  assign new_n5683_ = new_n9444_ & new_n9132_;
  assign new_n5684_ = new_n5683_ & new_n9113_;
  assign new_n5685_ = new_n9094_ & new_n9446_;
  assign new_n5686_ = new_n5685_ & new_n9151_;
  assign new_n5687_ = new_n9132_ & new_n9447_;
  assign new_n5688_ = new_n5687_ & new_n9151_;
  assign new_n5689_ = new_n5684_ | new_n5682_;
  assign new_n5690_ = new_n5689_ | new_n5686_;
  assign new_n5691_ = new_n5690_ | new_n5688_;
  assign new_n5692_ = new_n9409_ & new_n9239_;
  assign new_n5693_ = new_n5692_ & new_n9258_;
  assign new_n5694_ = new_n9413_ & new_n9277_;
  assign new_n5695_ = new_n5694_ & new_n9258_;
  assign new_n5696_ = new_n9239_ & new_n9448_;
  assign new_n5697_ = new_n5696_ & new_n9297_;
  assign new_n5698_ = new_n9277_ & new_n9449_;
  assign new_n5699_ = new_n5698_ & new_n9297_;
  assign new_n5700_ = new_n5695_ | new_n5693_;
  assign new_n5701_ = new_n5700_ | new_n5697_;
  assign new_n5702_ = new_n5701_ | new_n5699_;
  assign new_n5703_ = new_n5702_ & new_n9317_;
  assign new_n5704_ = new_n9439_ & new_n9241_;
  assign new_n5705_ = new_n5704_ & new_n9260_;
  assign new_n5706_ = new_n9443_ & new_n9279_;
  assign new_n5707_ = new_n5706_ & new_n9260_;
  assign new_n5708_ = new_n9241_ & new_n9450_;
  assign new_n5709_ = new_n5708_ & new_n9299_;
  assign new_n5710_ = new_n9279_ & new_n9451_;
  assign new_n5711_ = new_n5710_ & new_n9299_;
  assign new_n5712_ = new_n5707_ | new_n5705_;
  assign new_n5713_ = new_n5712_ | new_n5709_;
  assign new_n5714_ = new_n5713_ | new_n5711_;
  assign new_n5715_ = new_n5714_ & new_n9317_;
  assign new_n5716_ = new_n9429_ & new_n9242_;
  assign new_n5717_ = new_n5716_ & new_n9261_;
  assign new_n5718_ = new_n9433_ & new_n9280_;
  assign new_n5719_ = new_n5718_ & new_n9261_;
  assign new_n5720_ = new_n9242_ & new_n9452_;
  assign new_n5721_ = new_n5720_ & new_n9300_;
  assign new_n5722_ = new_n9280_ & new_n9453_;
  assign new_n5723_ = new_n5722_ & new_n9300_;
  assign new_n5724_ = new_n5719_ | new_n5717_;
  assign new_n5725_ = new_n5724_ | new_n5721_;
  assign new_n5726_ = new_n5725_ | new_n5723_;
  assign new_n5727_ = new_n5726_ & new_n9319_;
  assign new_n5728_ = new_n9419_ & new_n9244_;
  assign new_n5729_ = new_n5728_ & new_n9263_;
  assign new_n5730_ = new_n9423_ & new_n9282_;
  assign new_n5731_ = new_n5730_ & new_n9263_;
  assign new_n5732_ = new_n9244_ & new_n9454_;
  assign new_n5733_ = new_n5732_ & new_n9302_;
  assign new_n5734_ = new_n9282_ & new_n9455_;
  assign new_n5735_ = new_n5734_ & new_n9302_;
  assign new_n5736_ = new_n5731_ | new_n5729_;
  assign new_n5737_ = new_n5736_ | new_n5733_;
  assign new_n5738_ = new_n5737_ | new_n5735_;
  assign new_n5739_ = new_n5738_ & new_n9319_;
  assign new_n5740_ = new_n9411_ & new_n9337_;
  assign new_n5741_ = new_n5740_ & new_n9356_;
  assign new_n5742_ = new_n9415_ & new_n9375_;
  assign new_n5743_ = new_n5742_ & new_n9356_;
  assign new_n5744_ = new_n9337_ & new_n9448_;
  assign new_n5745_ = new_n5744_ & new_n9394_;
  assign new_n5746_ = new_n9375_ & new_n9449_;
  assign new_n5747_ = new_n5746_ & new_n9394_;
  assign new_n5748_ = new_n5743_ | new_n5741_;
  assign new_n5749_ = new_n5748_ | new_n5745_;
  assign new_n5750_ = new_n5749_ | new_n5747_;
  assign new_n5751_ = new_n5750_ & new_n9320_;
  assign new_n5752_ = new_n9441_ & new_n9339_;
  assign new_n5753_ = new_n5752_ & new_n9358_;
  assign new_n5754_ = new_n9445_ & new_n9377_;
  assign new_n5755_ = new_n5754_ & new_n9358_;
  assign new_n5756_ = new_n9339_ & new_n9450_;
  assign new_n5757_ = new_n5756_ & new_n9396_;
  assign new_n5758_ = new_n9377_ & new_n9451_;
  assign new_n5759_ = new_n5758_ & new_n9396_;
  assign new_n5760_ = new_n5755_ | new_n5753_;
  assign new_n5761_ = new_n5760_ | new_n5757_;
  assign new_n5762_ = new_n5761_ | new_n5759_;
  assign new_n5763_ = new_n5762_ & new_n9320_;
  assign new_n5764_ = new_n9431_ & new_n9340_;
  assign new_n5765_ = new_n5764_ & new_n9359_;
  assign new_n5766_ = new_n9435_ & new_n9378_;
  assign new_n5767_ = new_n5766_ & new_n9359_;
  assign new_n5768_ = new_n9340_ & new_n9452_;
  assign new_n5769_ = new_n5768_ & new_n9397_;
  assign new_n5770_ = new_n9378_ & new_n9453_;
  assign new_n5771_ = new_n5770_ & new_n9397_;
  assign new_n5772_ = new_n5767_ | new_n5765_;
  assign new_n5773_ = new_n5772_ | new_n5769_;
  assign new_n5774_ = new_n5773_ | new_n5771_;
  assign new_n5775_ = new_n5774_ & new_n9323_;
  assign new_n5776_ = new_n9421_ & new_n9342_;
  assign new_n5777_ = new_n5776_ & new_n9361_;
  assign new_n5778_ = new_n9425_ & new_n9380_;
  assign new_n5779_ = new_n5778_ & new_n9361_;
  assign new_n5780_ = new_n9342_ & new_n9454_;
  assign new_n5781_ = new_n5780_ & new_n9399_;
  assign new_n5782_ = new_n9380_ & new_n9455_;
  assign new_n5783_ = new_n5782_ & new_n9399_;
  assign new_n5784_ = new_n5779_ | new_n5777_;
  assign new_n5785_ = new_n5784_ | new_n5781_;
  assign new_n5786_ = new_n5785_ | new_n5783_;
  assign new_n5787_ = new_n5786_ & new_n9323_;
  assign new_n5788_ = new_n3823_ | new_n3179_;
  assign new_n5789_ = new_n9456_ & new_n9457_;
  assign new_n5790_ = new_n5789_ & new_n9458_;
  assign new_n5791_ = new_n9459_ & new_n9460_;
  assign new_n5792_ = new_n8789_ | new_n9461_;
  assign new_n5793_ = new_n9462_ & new_n9459_;
  assign new_n5794_ = new_n9463_ | new_n8789_;
  assign new_n5795_ = new_n9462_ & new_n9460_;
  assign new_n5796_ = new_n9463_ | new_n9461_;
  assign new_n5797_ = new_n5796_ & new_n5794_;
  assign new_n5798_ = new_n5795_ | new_n5793_;
  assign new_n5799_ = new_n9464_ & new_n9465_;
  assign new_n5800_ = new_n5799_ & new_n9458_;
  assign new_n5801_ = new_n9457_ & new_n9466_;
  assign new_n5802_ = new_n5801_ & new_n9467_;
  assign new_n5803_ = new_n9232_ & new_n9465_;
  assign new_n5804_ = new_n5803_ & new_n9467_;
  assign new_n5805_ = new_n5800_ | new_n5790_;
  assign new_n5806_ = new_n5805_ | new_n5802_;
  assign new_n5807_ = new_n5806_ | new_n5804_;
  assign new_n5808_ = new_n5807_ & new_n5788_;
  assign new_n5809_ = new_n5797_ | new_n9468_;
  assign new_n5810_ = new_n9469_ & new_n9464_;
  assign new_n5811_ = new_n9469_ & new_n9233_;
  assign new_n5812_ = new_n5811_ | new_n5810_;
  assign new_n5813_ = new_n9456_ & new_n8854_;
  assign new_n5814_ = new_n5813_ & new_n8894_;
  assign new_n5815_ = new_n9233_ & new_n8930_;
  assign new_n5816_ = new_n5815_ & new_n8896_;
  assign new_n5817_ = new_n8856_ & new_n9466_;
  assign new_n5818_ = new_n5817_ & new_n8953_;
  assign new_n5819_ = new_n5816_ | new_n5814_;
  assign new_n5820_ = new_n5819_ | new_n5818_;
  assign new_n5821_ = new_n8506_ & new_n8856_;
  assign new_n5822_ = new_n5821_ & new_n8896_;
  assign new_n5823_ = new_n9230_ & new_n8930_;
  assign new_n5824_ = new_n5823_ & new_n8897_;
  assign new_n5825_ = new_n8857_ & new_n3098_;
  assign new_n5826_ = new_n5825_ & new_n8953_;
  assign new_n5827_ = new_n5824_ | new_n5822_;
  assign new_n5828_ = new_n5827_ | new_n5826_;
  assign new_n5829_ = new_n8504_ & new_n8857_;
  assign new_n5830_ = new_n5829_ & new_n8897_;
  assign new_n5831_ = new_n9229_ & new_n8932_;
  assign new_n5832_ = new_n5831_ & new_n8901_;
  assign new_n5833_ = new_n8861_ & new_n3058_;
  assign new_n5834_ = new_n5833_ & new_n8955_;
  assign new_n5835_ = new_n5832_ | new_n5830_;
  assign new_n5836_ = new_n5835_ | new_n5834_;
  assign new_n5837_ = new_n8505_ & new_n8861_;
  assign new_n5838_ = new_n5837_ & new_n8901_;
  assign new_n5839_ = new_n9228_ & new_n8932_;
  assign new_n5840_ = new_n5839_ & new_n8902_;
  assign new_n5841_ = new_n8862_ & new_n3026_;
  assign new_n5842_ = new_n5841_ & new_n8955_;
  assign new_n5843_ = new_n5840_ | new_n5838_;
  assign new_n5844_ = new_n5843_ | new_n5842_;
  assign new_n5845_ = new_n9470_ | new_n8448_;
  assign new_n5846_ = new_n5845_ | new_n8447_;
  assign new_n5847_ = new_n5846_ | new_n9471_;
  assign new_n5848_ = new_n9472_ | new_n9473_;
  assign new_n5849_ = new_n5848_ | new_n9474_;
  assign new_n5850_ = new_n5849_ | new_n9475_;
  assign new_n5851_ = new_n5850_ | new_n9476_;
  assign new_n5852_ = new_n5851_ | new_n5847_;
  assign new_n5853_ = new_n5852_ | new_n9477_;
  assign new_n5854_ = new_n8831_ | new_n8782_;
  assign new_n5855_ = new_n5854_ | new_n9478_;
  assign new_n5856_ = new_n8832_ | new_n8781_;
  assign new_n5857_ = new_n5856_ | new_n9479_;
  assign new_n5858_ = new_n5857_ & new_n5855_;
  assign new_n5859_ = new_n3889_ & new_n9479_;
  assign new_n5860_ = new_n3891_ & new_n9478_;
  assign new_n5861_ = new_n5860_ | new_n5859_;
  assign new_n5862_ = new_n5861_ | new_n3572_;
  assign new_n5863_ = new_n5862_ & new_n5858_;
  assign new_n5864_ = new_n5863_ & new_n8862_;
  assign new_n5865_ = new_n5864_ & new_n8902_;
  assign new_n5866_ = new_n9227_ & new_n8933_;
  assign new_n5867_ = new_n5866_ & new_n8904_;
  assign new_n5868_ = new_n8864_ & new_n3050_;
  assign new_n5869_ = new_n5868_ & new_n8956_;
  assign new_n5870_ = new_n5867_ | new_n5865_;
  assign new_n5871_ = new_n5870_ | new_n5869_;
  assign new_n5872_ = new_n8581_ & new_n8864_;
  assign new_n5873_ = new_n5872_ & new_n8904_;
  assign new_n5874_ = new_n9226_ & new_n8933_;
  assign new_n5875_ = new_n5874_ & new_n8905_;
  assign new_n5876_ = new_n8865_ & new_n3042_;
  assign new_n5877_ = new_n5876_ & new_n8956_;
  assign new_n5878_ = new_n5875_ | new_n5873_;
  assign new_n5879_ = new_n5878_ | new_n5877_;
  assign new_n5880_ = new_n8580_ & new_n8865_;
  assign new_n5881_ = new_n5880_ & new_n8905_;
  assign new_n5882_ = new_n9225_ & new_n8936_;
  assign new_n5883_ = new_n5882_ & new_n8908_;
  assign new_n5884_ = new_n8868_ & new_n2842_;
  assign new_n5885_ = new_n5884_ & new_n8959_;
  assign new_n5886_ = new_n5883_ | new_n5881_;
  assign new_n5887_ = new_n5886_ | new_n5885_;
  assign new_n5888_ = new_n8578_ & new_n8868_;
  assign new_n5889_ = new_n5888_ & new_n8908_;
  assign new_n5890_ = new_n9224_ & new_n8936_;
  assign new_n5891_ = new_n5890_ & new_n8909_;
  assign new_n5892_ = new_n8869_ & new_n3034_;
  assign new_n5893_ = new_n5892_ & new_n8959_;
  assign new_n5894_ = new_n5891_ | new_n5889_;
  assign new_n5895_ = new_n5894_ | new_n5893_;
  assign new_n5896_ = new_n9482_ & new_n9095_;
  assign new_n5897_ = new_n5896_ & new_n9114_;
  assign new_n5898_ = new_n9486_ & new_n9133_;
  assign new_n5899_ = new_n5898_ & new_n9114_;
  assign new_n5900_ = new_n9095_ & new_n9488_;
  assign new_n5901_ = new_n5900_ & new_n9152_;
  assign new_n5902_ = new_n9133_ & new_n9489_;
  assign new_n5903_ = new_n5902_ & new_n9152_;
  assign new_n5904_ = new_n5899_ | new_n5897_;
  assign new_n5905_ = new_n5904_ | new_n5901_;
  assign new_n5906_ = new_n5905_ | new_n5903_;
  assign new_n5907_ = new_n9482_ & new_n9004_;
  assign new_n5908_ = new_n5907_ & new_n9023_;
  assign new_n5909_ = new_n9486_ & new_n9046_;
  assign new_n5910_ = new_n5909_ & new_n9023_;
  assign new_n5911_ = new_n9004_ & new_n9488_;
  assign new_n5912_ = new_n5911_ & new_n9066_;
  assign new_n5913_ = new_n9046_ & new_n9489_;
  assign new_n5914_ = new_n5913_ & new_n9066_;
  assign new_n5915_ = new_n5910_ | new_n5908_;
  assign new_n5916_ = new_n5915_ | new_n5912_;
  assign new_n5917_ = new_n5916_ | new_n5914_;
  assign new_n5918_ = new_n9492_ & new_n9007_;
  assign new_n5919_ = new_n5918_ & new_n9026_;
  assign new_n5920_ = new_n9496_ & new_n9049_;
  assign new_n5921_ = new_n5920_ & new_n9026_;
  assign new_n5922_ = new_n9007_ & new_n9498_;
  assign new_n5923_ = new_n5922_ & new_n9069_;
  assign new_n5924_ = new_n9049_ & new_n9499_;
  assign new_n5925_ = new_n5924_ & new_n9069_;
  assign new_n5926_ = new_n5921_ | new_n5919_;
  assign new_n5927_ = new_n5926_ | new_n5923_;
  assign new_n5928_ = new_n5927_ | new_n5925_;
  assign new_n5929_ = new_n9502_ & new_n9008_;
  assign new_n5930_ = new_n5929_ & new_n9027_;
  assign new_n5931_ = new_n9506_ & new_n9050_;
  assign new_n5932_ = new_n5931_ & new_n9027_;
  assign new_n5933_ = new_n9008_ & new_n9508_;
  assign new_n5934_ = new_n5933_ & new_n9070_;
  assign new_n5935_ = new_n9050_ & new_n9509_;
  assign new_n5936_ = new_n5935_ & new_n9070_;
  assign new_n5937_ = new_n5932_ | new_n5930_;
  assign new_n5938_ = new_n5937_ | new_n5934_;
  assign new_n5939_ = new_n5938_ | new_n5936_;
  assign new_n5940_ = new_n9512_ & new_n9010_;
  assign new_n5941_ = new_n5940_ & new_n9029_;
  assign new_n5942_ = new_n9516_ & new_n9052_;
  assign new_n5943_ = new_n5942_ & new_n9029_;
  assign new_n5944_ = new_n9010_ & new_n9518_;
  assign new_n5945_ = new_n5944_ & new_n9072_;
  assign new_n5946_ = new_n9052_ & new_n9519_;
  assign new_n5947_ = new_n5946_ & new_n9072_;
  assign new_n5948_ = new_n5943_ | new_n5941_;
  assign new_n5949_ = new_n5948_ | new_n5945_;
  assign new_n5950_ = new_n5949_ | new_n5947_;
  assign new_n5951_ = new_n9492_ & new_n9098_;
  assign new_n5952_ = new_n5951_ & new_n9117_;
  assign new_n5953_ = new_n9496_ & new_n9136_;
  assign new_n5954_ = new_n5953_ & new_n9117_;
  assign new_n5955_ = new_n9098_ & new_n9498_;
  assign new_n5956_ = new_n5955_ & new_n9155_;
  assign new_n5957_ = new_n9136_ & new_n9499_;
  assign new_n5958_ = new_n5957_ & new_n9155_;
  assign new_n5959_ = new_n5954_ | new_n5952_;
  assign new_n5960_ = new_n5959_ | new_n5956_;
  assign new_n5961_ = new_n5960_ | new_n5958_;
  assign new_n5962_ = new_n9502_ & new_n9099_;
  assign new_n5963_ = new_n5962_ & new_n9118_;
  assign new_n5964_ = new_n9506_ & new_n9137_;
  assign new_n5965_ = new_n5964_ & new_n9118_;
  assign new_n5966_ = new_n9099_ & new_n9508_;
  assign new_n5967_ = new_n5966_ & new_n9156_;
  assign new_n5968_ = new_n9137_ & new_n9509_;
  assign new_n5969_ = new_n5968_ & new_n9156_;
  assign new_n5970_ = new_n5965_ | new_n5963_;
  assign new_n5971_ = new_n5970_ | new_n5967_;
  assign new_n5972_ = new_n5971_ | new_n5969_;
  assign new_n5973_ = new_n9512_ & new_n9101_;
  assign new_n5974_ = new_n5973_ & new_n9120_;
  assign new_n5975_ = new_n9516_ & new_n9139_;
  assign new_n5976_ = new_n5975_ & new_n9120_;
  assign new_n5977_ = new_n9101_ & new_n9518_;
  assign new_n5978_ = new_n5977_ & new_n9158_;
  assign new_n5979_ = new_n9139_ & new_n9519_;
  assign new_n5980_ = new_n5979_ & new_n9158_;
  assign new_n5981_ = new_n5976_ | new_n5974_;
  assign new_n5982_ = new_n5981_ | new_n5978_;
  assign new_n5983_ = new_n5982_ | new_n5980_;
  assign new_n5984_ = new_n9511_ & new_n9245_;
  assign new_n5985_ = new_n5984_ & new_n9264_;
  assign new_n5986_ = new_n9515_ & new_n9283_;
  assign new_n5987_ = new_n5986_ & new_n9264_;
  assign new_n5988_ = new_n9245_ & new_n9520_;
  assign new_n5989_ = new_n5988_ & new_n9303_;
  assign new_n5990_ = new_n9283_ & new_n9521_;
  assign new_n5991_ = new_n5990_ & new_n9303_;
  assign new_n5992_ = new_n5987_ | new_n5985_;
  assign new_n5993_ = new_n5992_ | new_n5989_;
  assign new_n5994_ = new_n5993_ | new_n5991_;
  assign new_n5995_ = new_n5994_ & new_n9322_;
  assign new_n5996_ = new_n9501_ & new_n9248_;
  assign new_n5997_ = new_n5996_ & new_n9267_;
  assign new_n5998_ = new_n9505_ & new_n9286_;
  assign new_n5999_ = new_n5998_ & new_n9267_;
  assign new_n6000_ = new_n9248_ & new_n9522_;
  assign new_n6001_ = new_n6000_ & new_n9306_;
  assign new_n6002_ = new_n9286_ & new_n9523_;
  assign new_n6003_ = new_n6002_ & new_n9306_;
  assign new_n6004_ = new_n5999_ | new_n5997_;
  assign new_n6005_ = new_n6004_ | new_n6001_;
  assign new_n6006_ = new_n6005_ | new_n6003_;
  assign new_n6007_ = new_n6006_ & new_n9324_;
  assign new_n6008_ = new_n9491_ & new_n9249_;
  assign new_n6009_ = new_n6008_ & new_n9268_;
  assign new_n6010_ = new_n9495_ & new_n9287_;
  assign new_n6011_ = new_n6010_ & new_n9268_;
  assign new_n6012_ = new_n9249_ & new_n9524_;
  assign new_n6013_ = new_n6012_ & new_n9307_;
  assign new_n6014_ = new_n9287_ & new_n9525_;
  assign new_n6015_ = new_n6014_ & new_n9307_;
  assign new_n6016_ = new_n6011_ | new_n6009_;
  assign new_n6017_ = new_n6016_ | new_n6013_;
  assign new_n6018_ = new_n6017_ | new_n6015_;
  assign new_n6019_ = new_n6018_ & new_n9324_;
  assign new_n6020_ = new_n9481_ & new_n9251_;
  assign new_n6021_ = new_n6020_ & new_n9270_;
  assign new_n6022_ = new_n9485_ & new_n9289_;
  assign new_n6023_ = new_n6022_ & new_n9270_;
  assign new_n6024_ = new_n9251_ & new_n9526_;
  assign new_n6025_ = new_n6024_ & new_n9309_;
  assign new_n6026_ = new_n9289_ & new_n9527_;
  assign new_n6027_ = new_n6026_ & new_n9309_;
  assign new_n6028_ = new_n6023_ | new_n6021_;
  assign new_n6029_ = new_n6028_ | new_n6025_;
  assign new_n6030_ = new_n6029_ | new_n6027_;
  assign new_n6031_ = new_n6030_ & new_n9327_;
  assign new_n6032_ = new_n9513_ & new_n9343_;
  assign new_n6033_ = new_n6032_ & new_n9362_;
  assign new_n6034_ = new_n9517_ & new_n9381_;
  assign new_n6035_ = new_n6034_ & new_n9362_;
  assign new_n6036_ = new_n9343_ & new_n9520_;
  assign new_n6037_ = new_n6036_ & new_n9400_;
  assign new_n6038_ = new_n9381_ & new_n9521_;
  assign new_n6039_ = new_n6038_ & new_n9400_;
  assign new_n6040_ = new_n6035_ | new_n6033_;
  assign new_n6041_ = new_n6040_ | new_n6037_;
  assign new_n6042_ = new_n6041_ | new_n6039_;
  assign new_n6043_ = new_n6042_ & new_n9327_;
  assign new_n6044_ = new_n9503_ & new_n9346_;
  assign new_n6045_ = new_n6044_ & new_n9365_;
  assign new_n6046_ = new_n9507_ & new_n9384_;
  assign new_n6047_ = new_n6046_ & new_n9365_;
  assign new_n6048_ = new_n9346_ & new_n9522_;
  assign new_n6049_ = new_n6048_ & new_n9403_;
  assign new_n6050_ = new_n9384_ & new_n9523_;
  assign new_n6051_ = new_n6050_ & new_n9403_;
  assign new_n6052_ = new_n6047_ | new_n6045_;
  assign new_n6053_ = new_n6052_ | new_n6049_;
  assign new_n6054_ = new_n6053_ | new_n6051_;
  assign new_n6055_ = new_n6054_ & new_n9328_;
  assign new_n6056_ = new_n9493_ & new_n9347_;
  assign new_n6057_ = new_n6056_ & new_n9366_;
  assign new_n6058_ = new_n9497_ & new_n9385_;
  assign new_n6059_ = new_n6058_ & new_n9366_;
  assign new_n6060_ = new_n9347_ & new_n9524_;
  assign new_n6061_ = new_n6060_ & new_n9404_;
  assign new_n6062_ = new_n9385_ & new_n9525_;
  assign new_n6063_ = new_n6062_ & new_n9404_;
  assign new_n6064_ = new_n6059_ | new_n6057_;
  assign new_n6065_ = new_n6064_ | new_n6061_;
  assign new_n6066_ = new_n6065_ | new_n6063_;
  assign new_n6067_ = new_n6066_ & new_n9328_;
  assign new_n6068_ = new_n9483_ & new_n9349_;
  assign new_n6069_ = new_n6068_ & new_n9368_;
  assign new_n6070_ = new_n9487_ & new_n9387_;
  assign new_n6071_ = new_n6070_ & new_n9368_;
  assign new_n6072_ = new_n9349_ & new_n9526_;
  assign new_n6073_ = new_n6072_ & new_n9406_;
  assign new_n6074_ = new_n9387_ & new_n9527_;
  assign new_n6075_ = new_n6074_ & new_n9406_;
  assign new_n6076_ = new_n6071_ | new_n6069_;
  assign new_n6077_ = new_n6076_ | new_n6073_;
  assign new_n6078_ = new_n6077_ | new_n6075_;
  assign new_n6079_ = new_n6078_ & new_n9330_;
  assign new_n6080_ = new_n4449_ & new_n4435_;
  assign new_n6081_ = new_n4448_ & new_n4434_;
  assign new_n6082_ = new_n6081_ | new_n6080_;
  assign new_n6083_ = new_n9528_ | new_n8937_;
  assign new_n6084_ = new_n6083_ | new_n8960_;
  assign new_n6085_ = new_n4440_ | new_n4221_;
  assign new_n6086_ = new_n4442_ | new_n4219_;
  assign new_n6087_ = new_n6086_ & new_n6085_;
  assign new_n6088_ = new_n9529_ | new_n8869_;
  assign new_n6089_ = new_n6088_ | new_n8960_;
  assign new_n6090_ = new_n8937_ | new_n3091_;
  assign new_n6091_ = new_n6090_ | new_n8909_;
  assign new_n6092_ = new_n8911_ | new_n8871_;
  assign new_n6093_ = new_n6089_ & new_n6084_;
  assign new_n6094_ = new_n6093_ & new_n6091_;
  assign new_n6095_ = new_n6094_ & new_n9530_;
  assign new_n6096_ = new_n4446_ & new_n4433_;
  assign new_n6097_ = new_n4447_ & new_n4432_;
  assign new_n6098_ = new_n6097_ | new_n6096_;
  assign new_n6099_ = new_n9531_ | new_n8939_;
  assign new_n6100_ = new_n6099_ | new_n8962_;
  assign new_n6101_ = new_n4437_ | new_n4217_;
  assign new_n6102_ = new_n4438_ | new_n4214_;
  assign new_n6103_ = new_n6102_ & new_n6101_;
  assign new_n6104_ = new_n9532_ | new_n8871_;
  assign new_n6105_ = new_n6104_ | new_n8962_;
  assign new_n6106_ = new_n8939_ | new_n3075_;
  assign new_n6107_ = new_n6106_ | new_n8911_;
  assign new_n6108_ = new_n6105_ & new_n6100_;
  assign new_n6109_ = new_n6108_ & new_n6107_;
  assign new_n6110_ = new_n6109_ & new_n9530_;
  assign new_n6111_ = new_n9528_ & new_n8872_;
  assign new_n6112_ = new_n9529_ & new_n8940_;
  assign new_n6113_ = new_n6112_ | new_n6111_;
  assign new_n6114_ = new_n6113_ & new_n8912_;
  assign new_n6115_ = new_n8963_ & new_n2978_;
  assign new_n6116_ = new_n6115_ | new_n6114_;
  assign new_n6117_ = new_n9534_ & new_n9011_;
  assign new_n6118_ = new_n6117_ & new_n9030_;
  assign new_n6119_ = new_n9531_ & new_n8872_;
  assign new_n6120_ = new_n9532_ & new_n8940_;
  assign new_n6121_ = new_n6120_ | new_n6119_;
  assign new_n6122_ = new_n6121_ & new_n8912_;
  assign new_n6123_ = new_n8963_ & new_n2986_;
  assign new_n6124_ = new_n6123_ | new_n6122_;
  assign new_n6125_ = new_n9537_ & new_n9053_;
  assign new_n6126_ = new_n6125_ & new_n9030_;
  assign new_n6127_ = new_n9011_ & new_n9539_;
  assign new_n6128_ = new_n6127_ & new_n9073_;
  assign new_n6129_ = new_n9053_ & new_n9540_;
  assign new_n6130_ = new_n6129_ & new_n9073_;
  assign new_n6131_ = new_n6126_ | new_n6118_;
  assign new_n6132_ = new_n6131_ | new_n6128_;
  assign new_n6133_ = new_n6132_ | new_n6130_;
  assign new_n6134_ = new_n9534_ & new_n9102_;
  assign new_n6135_ = new_n6134_ & new_n9121_;
  assign new_n6136_ = new_n9537_ & new_n9140_;
  assign new_n6137_ = new_n6136_ & new_n9121_;
  assign new_n6138_ = new_n9102_ & new_n9539_;
  assign new_n6139_ = new_n6138_ & new_n9159_;
  assign new_n6140_ = new_n9140_ & new_n9540_;
  assign new_n6141_ = new_n6140_ & new_n9159_;
  assign new_n6142_ = new_n6137_ | new_n6135_;
  assign new_n6143_ = new_n6142_ | new_n6139_;
  assign new_n6144_ = new_n6143_ | new_n6141_;
  assign new_n6145_ = new_n9535_ & new_n9252_;
  assign new_n6146_ = new_n6145_ & new_n9271_;
  assign new_n6147_ = new_n9538_ & new_n9290_;
  assign new_n6148_ = new_n6147_ & new_n9271_;
  assign new_n6149_ = new_n9252_ & new_n9541_;
  assign new_n6150_ = new_n6149_ & new_n9310_;
  assign new_n6151_ = new_n9290_ & new_n9542_;
  assign new_n6152_ = new_n6151_ & new_n9310_;
  assign new_n6153_ = new_n6148_ | new_n6146_;
  assign new_n6154_ = new_n6153_ | new_n6150_;
  assign new_n6155_ = new_n6154_ | new_n6152_;
  assign new_n6156_ = new_n6155_ & new_n9330_;
  assign new_n6157_ = new_n9535_ & new_n9350_;
  assign new_n6158_ = new_n6157_ & new_n9369_;
  assign new_n6159_ = new_n9538_ & new_n9388_;
  assign new_n6160_ = new_n6159_ & new_n9369_;
  assign new_n6161_ = new_n9350_ & new_n9541_;
  assign new_n6162_ = new_n6161_ & new_n9407_;
  assign new_n6163_ = new_n9388_ & new_n9542_;
  assign new_n6164_ = new_n6163_ & new_n9407_;
  assign new_n6165_ = new_n6160_ | new_n6158_;
  assign new_n6166_ = new_n6165_ | new_n6162_;
  assign new_n6167_ = new_n6166_ | new_n6164_;
  assign new_n6168_ = new_n6167_ & new_n9331_;
  assign new_n6169_ = new_n4555_ & new_n4549_;
  assign new_n6170_ = new_n4554_ | new_n4548_;
  assign new_n6171_ = new_n9545_ & new_n9552_;
  assign new_n6172_ = new_n9557_ | new_n9563_;
  assign new_n6173_ = new_n6171_ & new_n4466_;
  assign new_n6174_ = new_n6172_ | new_n4467_;
  assign new_n6175_ = new_n9567_ & new_n9552_;
  assign new_n6176_ = new_n9573_ | new_n9563_;
  assign new_n6177_ = new_n6175_ & new_n4599_;
  assign new_n6178_ = new_n6176_ | new_n4598_;
  assign new_n6179_ = new_n6178_ & new_n6174_;
  assign new_n6180_ = new_n6177_ | new_n6173_;
  assign new_n6181_ = new_n9580_ & new_n9585_;
  assign new_n6182_ = new_n9589_ | new_n9594_;
  assign new_n6183_ = new_n9597_ & new_n9594_;
  assign new_n6184_ = new_n9603_ | new_n9585_;
  assign new_n6185_ = new_n6184_ & new_n6182_;
  assign new_n6186_ = new_n6183_ | new_n6181_;
  assign new_n6187_ = new_n6185_ & new_n9564_;
  assign new_n6188_ = new_n6186_ | new_n9551_;
  assign new_n6189_ = new_n6188_ & new_n6179_;
  assign new_n6190_ = new_n6187_ | new_n6180_;
  assign new_n6191_ = new_n3958_ & new_n9608_;
  assign new_n6192_ = new_n3959_ | new_n9609_;
  assign new_n6193_ = new_n6191_ & new_n9612_;
  assign new_n6194_ = new_n6192_ | new_n9618_;
  assign new_n6195_ = new_n6193_ & new_n9624_;
  assign new_n6196_ = new_n6194_ | new_n9629_;
  assign new_n6197_ = new_n6195_ & new_n9634_;
  assign new_n6198_ = new_n6196_ | new_n9638_;
  assign new_n6199_ = new_n3987_ & new_n9640_;
  assign new_n6200_ = new_n3986_ | new_n9641_;
  assign new_n6201_ = new_n6199_ & new_n9644_;
  assign new_n6202_ = new_n6200_ | new_n9650_;
  assign new_n6203_ = new_n6201_ & new_n9656_;
  assign new_n6204_ = new_n6202_ | new_n9661_;
  assign new_n6205_ = new_n6203_ & new_n9666_;
  assign new_n6206_ = new_n6204_ | new_n9670_;
  assign new_n6207_ = new_n9673_ & new_n9676_;
  assign new_n6208_ = new_n9679_ | new_n9681_;
  assign new_n6209_ = new_n9634_ & new_n4016_;
  assign new_n6210_ = new_n9638_ | new_n4017_;
  assign new_n6211_ = new_n9633_ & new_n9624_;
  assign new_n6212_ = new_n9637_ | new_n9629_;
  assign new_n6213_ = new_n6211_ & new_n3954_;
  assign new_n6214_ = new_n6212_ | new_n3955_;
  assign new_n6215_ = new_n9635_ & new_n9612_;
  assign new_n6216_ = new_n9639_ | new_n9618_;
  assign new_n6217_ = new_n6215_ & new_n3934_;
  assign new_n6218_ = new_n6216_ | new_n3935_;
  assign new_n6219_ = new_n6217_ & new_n9625_;
  assign new_n6220_ = new_n6218_ | new_n9630_;
  assign new_n6221_ = new_n9608_ & new_n9613_;
  assign new_n6222_ = new_n9609_ | new_n9619_;
  assign new_n6223_ = new_n6221_ & new_n9635_;
  assign new_n6224_ = new_n6222_ | new_n9639_;
  assign new_n6225_ = new_n6223_ & new_n3938_;
  assign new_n6226_ = new_n6224_ | new_n3939_;
  assign new_n6227_ = new_n6225_ & new_n9625_;
  assign new_n6228_ = new_n6226_ | new_n9630_;
  assign new_n6229_ = new_n6210_ & new_n6208_;
  assign new_n6230_ = new_n6209_ | new_n6207_;
  assign new_n6231_ = new_n6229_ & new_n6214_;
  assign new_n6232_ = new_n6230_ | new_n6213_;
  assign new_n6233_ = new_n6231_ & new_n6220_;
  assign new_n6234_ = new_n6232_ | new_n6219_;
  assign new_n6235_ = new_n6233_ & new_n6228_;
  assign new_n6236_ = new_n6234_ | new_n6227_;
  assign new_n6237_ = new_n9683_ & new_n9686_;
  assign new_n6238_ = new_n9689_ | new_n9691_;
  assign new_n6239_ = new_n9666_ & new_n4022_;
  assign new_n6240_ = new_n9670_ | new_n4023_;
  assign new_n6241_ = new_n9665_ & new_n9656_;
  assign new_n6242_ = new_n9669_ | new_n9661_;
  assign new_n6243_ = new_n6241_ & new_n3956_;
  assign new_n6244_ = new_n6242_ | new_n3957_;
  assign new_n6245_ = new_n9667_ & new_n9644_;
  assign new_n6246_ = new_n9671_ | new_n9650_;
  assign new_n6247_ = new_n6245_ & new_n3936_;
  assign new_n6248_ = new_n6246_ | new_n3937_;
  assign new_n6249_ = new_n6247_ & new_n9657_;
  assign new_n6250_ = new_n6248_ | new_n9662_;
  assign new_n6251_ = new_n9640_ & new_n9645_;
  assign new_n6252_ = new_n9641_ | new_n9651_;
  assign new_n6253_ = new_n6251_ & new_n9667_;
  assign new_n6254_ = new_n6252_ | new_n9671_;
  assign new_n6255_ = new_n6253_ & new_n3949_;
  assign new_n6256_ = new_n6254_ | new_n3948_;
  assign new_n6257_ = new_n6255_ & new_n9657_;
  assign new_n6258_ = new_n6256_ | new_n9662_;
  assign new_n6259_ = new_n6240_ & new_n6238_;
  assign new_n6260_ = new_n6239_ | new_n6237_;
  assign new_n6261_ = new_n6259_ & new_n6244_;
  assign new_n6262_ = new_n6260_ | new_n6243_;
  assign new_n6263_ = new_n6261_ & new_n6250_;
  assign new_n6264_ = new_n6262_ | new_n6249_;
  assign new_n6265_ = new_n6263_ & new_n6258_;
  assign new_n6266_ = new_n6264_ | new_n6257_;
  assign new_n6267_ = new_n9545_ & new_n9693_;
  assign new_n6268_ = new_n9557_ | new_n9695_;
  assign new_n6269_ = new_n9567_ & new_n9695_;
  assign new_n6270_ = new_n9573_ | new_n9693_;
  assign new_n6271_ = new_n6270_ & new_n6268_;
  assign new_n6272_ = new_n6269_ | new_n6267_;
  assign new_n6273_ = new_n4631_ & new_n4623_;
  assign new_n6274_ = new_n4630_ | new_n4622_;
  assign new_n6275_ = new_n4682_ & new_n4619_;
  assign new_n6276_ = new_n4683_ | new_n4618_;
  assign new_n6277_ = new_n4684_ & new_n4617_;
  assign new_n6278_ = new_n4685_ | new_n4616_;
  assign new_n6279_ = new_n6278_ & new_n6276_;
  assign new_n6280_ = new_n6277_ | new_n6275_;
  assign new_n6281_ = new_n9697_ & new_n9698_;
  assign new_n6282_ = new_n4483_ | new_n4481_;
  assign new_n6283_ = new_n9699_ & new_n9702_;
  assign new_n6284_ = new_n4135_ | new_n9704_;
  assign new_n6285_ = new_n9705_ & new_n3502_;
  assign new_n6286_ = new_n4098_ | new_n3503_;
  assign new_n6287_ = new_n6286_ & new_n6284_;
  assign new_n6288_ = new_n6285_ | new_n6283_;
  assign new_n6289_ = new_n9706_ & new_n9709_;
  assign new_n6290_ = new_n4137_ | new_n9711_;
  assign new_n6291_ = new_n9712_ & new_n3414_;
  assign new_n6292_ = new_n4100_ | new_n3415_;
  assign new_n6293_ = new_n6292_ & new_n6290_;
  assign new_n6294_ = new_n6291_ | new_n6289_;
  assign new_n6295_ = new_n9713_ & new_n9715_;
  assign new_n6296_ = new_n4689_ | new_n9716_;
  assign new_n6297_ = new_n9717_ & new_n9718_;
  assign new_n6298_ = new_n4691_ | new_n9720_;
  assign new_n6299_ = new_n6298_ & new_n6296_;
  assign new_n6300_ = new_n6297_ | new_n6295_;
  assign new_n6301_ = new_n9722_ & new_n9726_;
  assign new_n6302_ = new_n9731_ & new_n9734_;
  assign new_n6303_ = new_n9738_ | new_n9741_;
  assign new_n6304_ = new_n9744_ | new_n9747_;
  assign new_n6305_ = new_n9749_ & new_n9750_;
  assign new_n6306_ = new_n4677_ | new_n4673_;
  assign new_n6307_ = new_n9751_ & new_n9752_;
  assign new_n6308_ = new_n4681_ | new_n4669_;
  assign new_n6309_ = new_n9754_ & new_n9756_;
  assign new_n6310_ = new_n9758_ & new_n9761_;
  assign new_n6311_ = new_n6310_ | new_n6309_;
  assign new_n6312_ = new_n9731_ & new_n9765_;
  assign new_n6313_ = new_n9767_ & new_n9734_;
  assign new_n6314_ = new_n6313_ | new_n6312_;
  assign new_n6315_ = new_n9769_ & new_n9741_;
  assign new_n6316_ = new_n9738_ | new_n9773_;
  assign new_n6317_ = new_n9737_ & new_n9773_;
  assign new_n6318_ = new_n9769_ | new_n9742_;
  assign new_n6319_ = new_n6318_ & new_n6316_;
  assign new_n6320_ = new_n6317_ | new_n6315_;
  assign new_n6321_ = new_n9778_ & new_n9782_;
  assign new_n6322_ = new_n9785_ | new_n9788_;
  assign new_n6323_ = new_n9790_ & new_n9791_;
  assign new_n6324_ = new_n9792_ | new_n9793_;
  assign new_n6325_ = new_n9792_ & new_n9793_;
  assign new_n6326_ = new_n9790_ | new_n9791_;
  assign new_n6327_ = new_n6326_ & new_n6324_;
  assign new_n6328_ = new_n6325_ | new_n6323_;
  assign new_n6329_ = new_n9794_ & new_n9795_;
  assign new_n6330_ = new_n9796_ | new_n9797_;
  assign new_n6331_ = new_n9796_ & new_n9797_;
  assign new_n6332_ = new_n9794_ | new_n9795_;
  assign new_n6333_ = new_n6332_ & new_n6330_;
  assign new_n6334_ = new_n6331_ | new_n6329_;
  assign new_n6335_ = new_n9798_ & new_n9799_;
  assign new_n6336_ = new_n9800_ | new_n9801_;
  assign new_n6337_ = new_n9800_ & new_n9801_;
  assign new_n6338_ = new_n9798_ | new_n9799_;
  assign new_n6339_ = new_n6338_ & new_n6336_;
  assign new_n6340_ = new_n6337_ | new_n6335_;
  assign new_n6341_ = new_n9802_ & new_n9803_;
  assign new_n6342_ = new_n9804_ | new_n9805_;
  assign new_n6343_ = new_n9804_ & new_n9805_;
  assign new_n6344_ = new_n9802_ | new_n9803_;
  assign new_n6345_ = new_n6344_ & new_n6342_;
  assign new_n6346_ = new_n6343_ | new_n6341_;
  assign new_n6347_ = new_n9806_ & new_n9807_;
  assign new_n6348_ = new_n4675_ | new_n4671_;
  assign new_n6349_ = new_n9808_ & new_n9809_;
  assign new_n6350_ = new_n4679_ | new_n4667_;
  assign new_n6351_ = new_n9778_ & new_n9788_;
  assign new_n6352_ = new_n9785_ | new_n9782_;
  assign new_n6353_ = new_n9786_ & new_n9781_;
  assign new_n6354_ = new_n9777_ | new_n9789_;
  assign new_n6355_ = new_n6354_ & new_n6352_;
  assign new_n6356_ = new_n6353_ | new_n6351_;
  assign new_n6357_ = new_n9718_ & new_n9810_;
  assign new_n6358_ = new_n9720_ | new_n3505_;
  assign new_n6359_ = new_n6358_ & new_n9716_;
  assign new_n6360_ = new_n6357_ | new_n9715_;
  assign new_n6361_ = new_n9811_ & new_n9812_;
  assign new_n6362_ = new_n4507_ | new_n3441_;
  assign new_n6363_ = new_n4259_ & new_n3444_;
  assign new_n6364_ = new_n9813_ | new_n3445_;
  assign new_n6365_ = new_n6364_ & new_n6362_;
  assign new_n6366_ = new_n6363_ | new_n6361_;
  assign new_n6367_ = new_n9816_ & new_n9820_;
  assign new_n6368_ = new_n9823_ | new_n3483_;
  assign new_n6369_ = new_n9823_ & new_n3486_;
  assign new_n6370_ = new_n9816_ | new_n3487_;
  assign new_n6371_ = new_n6370_ & new_n6368_;
  assign new_n6372_ = new_n6369_ | new_n6367_;
  assign new_n6373_ = new_n9827_ & new_n9831_;
  assign new_n6374_ = new_n9834_ | new_n3395_;
  assign new_n6375_ = new_n9834_ & new_n3398_;
  assign new_n6376_ = new_n9827_ | new_n3399_;
  assign new_n6377_ = new_n6376_ & new_n6374_;
  assign new_n6378_ = new_n6375_ | new_n6373_;
  assign new_n6379_ = new_n9754_ & new_n9761_;
  assign new_n6380_ = new_n4607_ & new_n4297_;
  assign new_n6381_ = new_n4606_ | new_n4296_;
  assign new_n6382_ = new_n4584_ & new_n4474_;
  assign new_n6383_ = new_n4585_ | new_n4475_;
  assign new_n6384_ = new_n6383_ & new_n6381_;
  assign new_n6385_ = new_n6382_ | new_n6380_;
  assign new_n6386_ = new_n9836_ & new_n9838_;
  assign new_n6387_ = new_n9840_ | new_n9843_;
  assign new_n6388_ = new_n9840_ & new_n9843_;
  assign new_n6389_ = new_n9836_ | new_n9838_;
  assign new_n6390_ = new_n6389_ & new_n6387_;
  assign new_n6391_ = new_n6388_ | new_n6386_;
  assign new_n6392_ = new_n6391_ | new_n9846_;
  assign new_n6393_ = new_n6390_ | new_n9847_;
  assign new_n6394_ = new_n6393_ & new_n6392_;
  assign new_n6395_ = new_n9848_ | new_n9850_;
  assign new_n6396_ = new_n6395_ | new_n9852_;
  assign new_n6397_ = new_n4605_ & new_n4295_;
  assign new_n6398_ = new_n4604_ | new_n4294_;
  assign new_n6399_ = new_n4582_ & new_n4472_;
  assign new_n6400_ = new_n4583_ | new_n4473_;
  assign new_n6401_ = new_n6400_ & new_n6398_;
  assign new_n6402_ = new_n6399_ | new_n6397_;
  assign new_n6403_ = new_n9853_ & new_n9839_;
  assign new_n6404_ = new_n9854_ | new_n9842_;
  assign new_n6405_ = new_n9854_ & new_n9844_;
  assign new_n6406_ = new_n9853_ | new_n9839_;
  assign new_n6407_ = new_n6406_ & new_n6404_;
  assign new_n6408_ = new_n6405_ | new_n6403_;
  assign new_n6409_ = new_n6408_ | new_n9846_;
  assign new_n6410_ = new_n6407_ | new_n9847_;
  assign new_n6411_ = new_n6410_ & new_n6409_;
  assign new_n6412_ = new_n9855_ | new_n9856_;
  assign new_n6413_ = new_n6412_ | new_n9852_;
  assign new_n6414_ = new_n9856_ & new_n6198_;
  assign new_n6415_ = new_n9850_ | new_n9857_;
  assign new_n6416_ = new_n6415_ | new_n9848_;
  assign new_n6417_ = new_n6416_ | new_n9859_;
  assign new_n6418_ = new_n6414_ | new_n9855_;
  assign new_n6419_ = new_n6418_ | new_n9859_;
  assign new_n6420_ = new_n6413_ & new_n6396_;
  assign new_n6421_ = new_n6420_ & new_n6417_;
  assign new_n6422_ = new_n6421_ & new_n6419_;
  assign new_n6423_ = new_n4556_ & new_n4551_;
  assign new_n6424_ = new_n4557_ | new_n4550_;
  assign new_n6425_ = new_n9860_ & new_n9619_;
  assign new_n6426_ = new_n9861_ | new_n9613_;
  assign new_n6427_ = new_n9861_ & new_n9615_;
  assign new_n6428_ = new_n9860_ | new_n9621_;
  assign new_n6429_ = new_n6428_ & new_n6426_;
  assign new_n6430_ = new_n6427_ | new_n6425_;
  assign new_n6431_ = new_n6430_ | new_n9626_;
  assign new_n6432_ = new_n6429_ | new_n9631_;
  assign new_n6433_ = new_n6432_ & new_n6431_;
  assign new_n6434_ = new_n6433_ & new_n9858_;
  assign new_n6435_ = new_n4600_ & new_n4451_;
  assign new_n6436_ = new_n4601_ | new_n4450_;
  assign new_n6437_ = new_n4594_ & new_n4469_;
  assign new_n6438_ = new_n4595_ | new_n4468_;
  assign new_n6439_ = new_n6438_ & new_n6436_;
  assign new_n6440_ = new_n6437_ | new_n6435_;
  assign new_n6441_ = new_n9862_ & new_n9621_;
  assign new_n6442_ = new_n9863_ | new_n9615_;
  assign new_n6443_ = new_n9863_ & new_n9614_;
  assign new_n6444_ = new_n9862_ | new_n9620_;
  assign new_n6445_ = new_n6444_ & new_n6442_;
  assign new_n6446_ = new_n6443_ | new_n6441_;
  assign new_n6447_ = new_n6445_ & new_n9631_;
  assign new_n6448_ = new_n6446_ & new_n9626_;
  assign new_n6449_ = new_n6448_ | new_n6447_;
  assign new_n6450_ = new_n6449_ & new_n9851_;
  assign new_n6451_ = new_n6450_ | new_n6434_;
  assign new_n6452_ = new_n4610_ & new_n4301_;
  assign new_n6453_ = new_n4611_ | new_n4300_;
  assign new_n6454_ = new_n4588_ & new_n4479_;
  assign new_n6455_ = new_n4589_ | new_n4478_;
  assign new_n6456_ = new_n6455_ & new_n6453_;
  assign new_n6457_ = new_n6454_ | new_n6452_;
  assign new_n6458_ = new_n9864_ & new_n9868_;
  assign new_n6459_ = new_n9874_ | new_n9876_;
  assign new_n6460_ = new_n9874_ & new_n9876_;
  assign new_n6461_ = new_n9864_ | new_n9868_;
  assign new_n6462_ = new_n6461_ & new_n6459_;
  assign new_n6463_ = new_n6460_ | new_n6458_;
  assign new_n6464_ = new_n6462_ & new_n9879_;
  assign new_n6465_ = new_n6463_ & new_n9880_;
  assign new_n6466_ = new_n6465_ | new_n6464_;
  assign new_n6467_ = new_n9881_ & new_n9882_;
  assign new_n6468_ = new_n6467_ & new_n9884_;
  assign new_n6469_ = new_n4608_ & new_n4299_;
  assign new_n6470_ = new_n4609_ | new_n4298_;
  assign new_n6471_ = new_n4586_ & new_n4477_;
  assign new_n6472_ = new_n4587_ | new_n4476_;
  assign new_n6473_ = new_n6472_ & new_n6470_;
  assign new_n6474_ = new_n6471_ | new_n6469_;
  assign new_n6475_ = new_n9885_ & new_n9869_;
  assign new_n6476_ = new_n9886_ | new_n9877_;
  assign new_n6477_ = new_n9886_ & new_n9877_;
  assign new_n6478_ = new_n9885_ | new_n9869_;
  assign new_n6479_ = new_n6478_ & new_n6476_;
  assign new_n6480_ = new_n6477_ | new_n6475_;
  assign new_n6481_ = new_n6479_ & new_n9879_;
  assign new_n6482_ = new_n6480_ & new_n9880_;
  assign new_n6483_ = new_n6482_ | new_n6481_;
  assign new_n6484_ = new_n9887_ & new_n9889_;
  assign new_n6485_ = new_n6484_ & new_n9884_;
  assign new_n6486_ = new_n9882_ & new_n6206_;
  assign new_n6487_ = new_n9889_ | new_n9890_;
  assign new_n6488_ = new_n6486_ & new_n9881_;
  assign new_n6489_ = new_n6488_ & new_n9892_;
  assign new_n6490_ = new_n6487_ & new_n9887_;
  assign new_n6491_ = new_n6490_ & new_n9892_;
  assign new_n6492_ = new_n6485_ | new_n6468_;
  assign new_n6493_ = new_n6492_ | new_n6489_;
  assign new_n6494_ = new_n6493_ | new_n6491_;
  assign new_n6495_ = new_n4558_ & new_n4553_;
  assign new_n6496_ = new_n4559_ | new_n4552_;
  assign new_n6497_ = new_n9893_ & new_n9651_;
  assign new_n6498_ = new_n9894_ | new_n9645_;
  assign new_n6499_ = new_n9894_ & new_n9647_;
  assign new_n6500_ = new_n9893_ | new_n9653_;
  assign new_n6501_ = new_n6500_ & new_n6498_;
  assign new_n6502_ = new_n6499_ | new_n6497_;
  assign new_n6503_ = new_n6502_ | new_n9658_;
  assign new_n6504_ = new_n6501_ | new_n9663_;
  assign new_n6505_ = new_n6504_ & new_n6503_;
  assign new_n6506_ = new_n6505_ & new_n9883_;
  assign new_n6507_ = new_n4602_ & new_n4453_;
  assign new_n6508_ = new_n4603_ | new_n4452_;
  assign new_n6509_ = new_n4596_ & new_n4471_;
  assign new_n6510_ = new_n4597_ | new_n4470_;
  assign new_n6511_ = new_n6510_ & new_n6508_;
  assign new_n6512_ = new_n6509_ | new_n6507_;
  assign new_n6513_ = new_n9895_ & new_n9653_;
  assign new_n6514_ = new_n9896_ | new_n9647_;
  assign new_n6515_ = new_n9896_ & new_n9646_;
  assign new_n6516_ = new_n9895_ | new_n9652_;
  assign new_n6517_ = new_n6516_ & new_n6514_;
  assign new_n6518_ = new_n6515_ | new_n6513_;
  assign new_n6519_ = new_n6517_ & new_n9663_;
  assign new_n6520_ = new_n6518_ & new_n9658_;
  assign new_n6521_ = new_n6520_ | new_n6519_;
  assign new_n6522_ = new_n6521_ & new_n9891_;
  assign new_n6523_ = new_n6522_ | new_n6506_;
  assign new_n6524_ = new_n9722_ & new_n9898_;
  assign new_n6525_ = new_n9900_ & new_n9726_;
  assign new_n6526_ = new_n6525_ | new_n6524_;
  assign new_n6527_ = new_n9902_ & new_n9564_;
  assign new_n6528_ = new_n9903_ & new_n9553_;
  assign new_n6529_ = new_n6528_ | new_n6527_;
  assign new_n6530_ = new_n9905_ & new_n9747_;
  assign new_n6531_ = new_n9744_ & new_n9909_;
  assign new_n6532_ = new_n6531_ | new_n6530_;
  assign new_n6533_ = new_n9706_ & new_n9914_;
  assign new_n6534_ = new_n9712_ & new_n3386_;
  assign new_n6535_ = new_n6534_ | new_n6533_;
  assign new_n6536_ = new_n6293_ & new_n9917_;
  assign new_n6537_ = new_n9919_ & new_n3565_;
  assign new_n6538_ = new_n6537_ | new_n6536_;
  assign new_n6539_ = new_n6287_ & new_n9921_;
  assign new_n6540_ = new_n9923_ & new_n3593_;
  assign new_n6541_ = new_n6540_ | new_n6539_;
  assign new_n6542_ = new_n9817_ & new_n9924_;
  assign new_n6543_ = new_n9822_ | new_n3489_;
  assign new_n6544_ = new_n9824_ & new_n3492_;
  assign new_n6545_ = new_n9817_ | new_n3493_;
  assign new_n6546_ = new_n6545_ & new_n6543_;
  assign new_n6547_ = new_n6544_ | new_n6542_;
  assign new_n6548_ = new_n9828_ & new_n9925_;
  assign new_n6549_ = new_n9833_ | new_n3401_;
  assign new_n6550_ = new_n9835_ & new_n3404_;
  assign new_n6551_ = new_n9828_ | new_n3405_;
  assign new_n6552_ = new_n6551_ & new_n6549_;
  assign new_n6553_ = new_n6550_ | new_n6548_;
  assign new_n6554_ = new_n9927_ & new_n9931_;
  assign new_n6555_ = new_n9935_ & new_n9938_;
  assign new_n6556_ = new_n9941_ & new_n9945_;
  assign new_n6557_ = new_n9949_ & new_n9953_;
  assign new_n6558_ = new_n9723_ | new_n9727_;
  assign new_n6559_ = new_n9905_ | new_n9909_;
  assign new_n6560_ = new_n9957_ & new_n9960_;
  assign new_n6561_ = new_n9963_ & new_n9966_;
  assign new_n6562_ = new_n9970_ & new_n9973_;
  assign new_n6563_ = new_n9976_ & new_n3869_;
  assign new_n6564_ = new_n3871_ & new_n9977_;
  assign new_n6565_ = new_n9980_ & new_n9982_;
  assign new_n6566_ = new_n9985_ & new_n9988_;
  assign new_n6567_ = new_n9989_ & new_n3873_;
  assign new_n6568_ = new_n3877_ & new_n9990_;
  assign new_n6569_ = new_n9692_ & new_n9991_;
  assign new_n6570_ = new_n9696_ & new_n3525_;
  assign new_n6571_ = new_n9993_ & new_n9995_;
  assign new_n6572_ = new_n9997_ & new_n10000_;
  assign new_n6573_ = new_n10000_ & new_n10003_;
  assign new_n6574_ = new_n9997_ | new_n10003_;
  assign new_n6575_ = new_n10005_ | new_n10008_;
  assign new_n6576_ = new_n6319_ | new_n10013_;
  assign new_n6577_ = new_n10015_ & new_n10005_;
  assign new_n6578_ = new_n10015_ | new_n10008_;
  assign new_n6579_ = new_n9970_ & new_n10016_;
  assign new_n6580_ = new_n10017_ & new_n9963_;
  assign new_n6581_ = new_n3880_ & new_n9991_;
  assign new_n6582_ = new_n3857_ & new_n3530_;
  assign new_n6583_ = new_n6582_ | new_n6581_;
  assign new_n6584_ = new_n10018_ | new_n10020_;
  assign new_n6585_ = new_n9753_ & new_n9767_;
  assign new_n6586_ = new_n9673_ & new_n9900_;
  assign new_n6587_ = new_n9758_ & new_n9730_;
  assign new_n6588_ = new_n10022_ & new_n10024_;
  assign new_n6589_ = new_n10025_ & new_n4031_;
  assign new_n6590_ = new_n9679_ & new_n9723_;
  assign new_n6591_ = new_n10018_ & new_n10020_;
  assign new_n6592_ = new_n10026_ & new_n9993_;
  assign new_n6593_ = new_n10027_ & new_n9999_;
  assign new_n6594_ = new_n10028_ | new_n10029_;
  assign new_n6595_ = new_n6594_ | new_n10030_;
  assign new_n6596_ = new_n10031_ & new_n10009_;
  assign new_n6597_ = new_n6596_ & new_n10032_;
  assign new_n6598_ = new_n10033_ & new_n3929_;
  assign new_n6599_ = new_n4037_ & new_n10034_;
  assign new_n6600_ = new_n6599_ | new_n6598_;
  assign new_n6601_ = new_n9927_ & new_n10036_;
  assign new_n6602_ = new_n3919_ & new_n9931_;
  assign new_n6603_ = new_n6602_ | new_n6601_;
  assign new_n6604_ = new_n9935_ & new_n10038_;
  assign new_n6605_ = new_n3971_ & new_n9938_;
  assign new_n6606_ = new_n6605_ | new_n6604_;
  assign new_n6607_ = new_n9941_ & new_n10040_;
  assign new_n6608_ = new_n3909_ & new_n9945_;
  assign new_n6609_ = new_n6608_ | new_n6607_;
  assign new_n6610_ = new_n9949_ & new_n10043_;
  assign new_n6611_ = new_n3911_ & new_n9953_;
  assign new_n6612_ = new_n6611_ | new_n6610_;
  assign new_n6613_ = new_n9674_ & new_n9681_;
  assign new_n6614_ = new_n9678_ & new_n9676_;
  assign new_n6615_ = new_n6614_ | new_n6613_;
  assign new_n6616_ = new_n9683_ & new_n9691_;
  assign new_n6617_ = new_n9689_ & new_n9686_;
  assign new_n6618_ = new_n6617_ | new_n6616_;
  assign new_n6619_ = new_n9957_ & new_n10046_;
  assign new_n6620_ = new_n10047_ & new_n9960_;
  assign new_n6621_ = new_n6620_ | new_n6619_;
  assign new_n6622_ = new_n9962_ & new_n10049_;
  assign new_n6623_ = new_n10016_ & new_n9966_;
  assign new_n6624_ = new_n6623_ | new_n6622_;
  assign new_n6625_ = new_n9969_ & new_n10052_;
  assign new_n6626_ = new_n10017_ & new_n9973_;
  assign new_n6627_ = new_n6626_ | new_n6625_;
  assign new_n6628_ = new_n9684_ & new_n10047_;
  assign new_n6629_ = new_n9688_ & new_n9956_;
  assign new_n6630_ = new_n6629_ | new_n6628_;
  assign new_n6631_ = new_n3882_ & new_n9982_;
  assign new_n6632_ = new_n3883_ | new_n9988_;
  assign new_n6633_ = new_n3859_ & new_n3462_;
  assign new_n6634_ = new_n3858_ | new_n3463_;
  assign new_n6635_ = new_n6634_ & new_n6632_;
  assign new_n6636_ = new_n6633_ | new_n6631_;
  assign new_n6637_ = new_n6636_ | new_n9902_;
  assign new_n6638_ = new_n6635_ | new_n9903_;
  assign new_n6639_ = new_n6638_ & new_n6637_;
  assign new_n6640_ = new_n10056_ & new_n9727_;
  assign new_n6641_ = new_n10061_ | new_n9898_;
  assign new_n6642_ = new_n6640_ & new_n10065_;
  assign new_n6643_ = new_n6641_ | new_n10066_;
  assign new_n6644_ = new_n10069_ & new_n9729_;
  assign new_n6645_ = new_n10074_ | new_n9899_;
  assign new_n6646_ = new_n6644_ & new_n10066_;
  assign new_n6647_ = new_n6645_ | new_n10065_;
  assign new_n6648_ = new_n6647_ & new_n6643_;
  assign new_n6649_ = new_n6646_ | new_n6642_;
  assign new_n6650_ = new_n10080_ & new_n10085_;
  assign new_n6651_ = new_n10089_ | new_n10096_;
  assign new_n6652_ = new_n10100_ & new_n10096_;
  assign new_n6653_ = new_n10108_ | new_n10085_;
  assign new_n6654_ = new_n6653_ & new_n6651_;
  assign new_n6655_ = new_n6652_ | new_n6650_;
  assign new_n6656_ = new_n6654_ & new_n9899_;
  assign new_n6657_ = new_n6655_ | new_n9729_;
  assign new_n6658_ = new_n6657_ & new_n6648_;
  assign new_n6659_ = new_n6656_ | new_n6649_;
  assign new_n6660_ = new_n10056_ & new_n9735_;
  assign new_n6661_ = new_n10061_ | new_n9765_;
  assign new_n6662_ = new_n6660_ & new_n10113_;
  assign new_n6663_ = new_n6661_ | new_n10114_;
  assign new_n6664_ = new_n10069_ & new_n9735_;
  assign new_n6665_ = new_n10074_ | new_n9766_;
  assign new_n6666_ = new_n6664_ & new_n10114_;
  assign new_n6667_ = new_n6665_ | new_n10113_;
  assign new_n6668_ = new_n6667_ & new_n6663_;
  assign new_n6669_ = new_n6666_ | new_n6662_;
  assign new_n6670_ = new_n10080_ & new_n10115_;
  assign new_n6671_ = new_n10089_ | new_n10118_;
  assign new_n6672_ = new_n10100_ & new_n10118_;
  assign new_n6673_ = new_n10108_ | new_n10115_;
  assign new_n6674_ = new_n6673_ & new_n6671_;
  assign new_n6675_ = new_n6672_ | new_n6670_;
  assign new_n6676_ = new_n6674_ & new_n9766_;
  assign new_n6677_ = new_n6675_ | new_n9736_;
  assign new_n6678_ = new_n6677_ & new_n6668_;
  assign new_n6679_ = new_n6676_ | new_n6669_;
  assign new_n6680_ = new_n10120_ & new_n10121_;
  assign new_n6681_ = new_n10122_ | new_n10123_;
  assign new_n6682_ = new_n10122_ & new_n10123_;
  assign new_n6683_ = new_n10120_ | new_n10121_;
  assign new_n6684_ = new_n6683_ & new_n6681_;
  assign new_n6685_ = new_n6682_ | new_n6680_;
  assign new_n6686_ = new_n10057_ & new_n9762_;
  assign new_n6687_ = new_n10062_ | new_n9756_;
  assign new_n6688_ = new_n6686_ & new_n10124_;
  assign new_n6689_ = new_n6687_ | new_n10125_;
  assign new_n6690_ = new_n10070_ & new_n9762_;
  assign new_n6691_ = new_n10075_ | new_n9757_;
  assign new_n6692_ = new_n6690_ & new_n10125_;
  assign new_n6693_ = new_n6691_ | new_n10124_;
  assign new_n6694_ = new_n6693_ & new_n6689_;
  assign new_n6695_ = new_n6692_ | new_n6688_;
  assign new_n6696_ = new_n10081_ & new_n10126_;
  assign new_n6697_ = new_n10088_ | new_n10129_;
  assign new_n6698_ = new_n10101_ & new_n10129_;
  assign new_n6699_ = new_n10107_ | new_n10126_;
  assign new_n6700_ = new_n6699_ & new_n6697_;
  assign new_n6701_ = new_n6698_ | new_n6696_;
  assign new_n6702_ = new_n6700_ & new_n9757_;
  assign new_n6703_ = new_n6701_ | new_n9763_;
  assign new_n6704_ = new_n6703_ & new_n6694_;
  assign new_n6705_ = new_n6702_ | new_n6695_;
  assign new_n6706_ = new_n10131_ & new_n10132_;
  assign new_n6707_ = new_n10133_ | new_n10135_;
  assign new_n6708_ = new_n10133_ & new_n10135_;
  assign new_n6709_ = new_n10131_ | new_n10132_;
  assign new_n6710_ = new_n6709_ & new_n6707_;
  assign new_n6711_ = new_n6708_ | new_n6706_;
  assign new_n6712_ = new_n6711_ | new_n6684_;
  assign new_n6713_ = new_n6710_ | new_n6685_;
  assign new_n6714_ = new_n6713_ & new_n6712_;
  assign new_n6715_ = new_n9546_ & new_n9910_;
  assign new_n6716_ = new_n9556_ | new_n9746_;
  assign new_n6717_ = new_n6715_ & new_n10136_;
  assign new_n6718_ = new_n6716_ | new_n10137_;
  assign new_n6719_ = new_n9568_ & new_n9910_;
  assign new_n6720_ = new_n9574_ | new_n9748_;
  assign new_n6721_ = new_n6719_ & new_n10137_;
  assign new_n6722_ = new_n6720_ | new_n10136_;
  assign new_n6723_ = new_n6722_ & new_n6718_;
  assign new_n6724_ = new_n6721_ | new_n6717_;
  assign new_n6725_ = new_n9580_ & new_n10138_;
  assign new_n6726_ = new_n9589_ | new_n10141_;
  assign new_n6727_ = new_n9597_ & new_n10141_;
  assign new_n6728_ = new_n9603_ | new_n10138_;
  assign new_n6729_ = new_n6728_ & new_n6726_;
  assign new_n6730_ = new_n6727_ | new_n6725_;
  assign new_n6731_ = new_n6729_ & new_n9748_;
  assign new_n6732_ = new_n6730_ | new_n9911_;
  assign new_n6733_ = new_n6732_ & new_n6723_;
  assign new_n6734_ = new_n6731_ | new_n6724_;
  assign new_n6735_ = new_n9546_ & new_n9774_;
  assign new_n6736_ = new_n9558_ | new_n9742_;
  assign new_n6737_ = new_n6735_ & new_n10143_;
  assign new_n6738_ = new_n6736_ | new_n10144_;
  assign new_n6739_ = new_n9568_ & new_n9774_;
  assign new_n6740_ = new_n9574_ | new_n9743_;
  assign new_n6741_ = new_n6739_ & new_n10144_;
  assign new_n6742_ = new_n6740_ | new_n10143_;
  assign new_n6743_ = new_n6742_ & new_n6738_;
  assign new_n6744_ = new_n6741_ | new_n6737_;
  assign new_n6745_ = new_n9581_ & new_n10145_;
  assign new_n6746_ = new_n9588_ | new_n10148_;
  assign new_n6747_ = new_n9598_ & new_n10148_;
  assign new_n6748_ = new_n9604_ | new_n10145_;
  assign new_n6749_ = new_n6748_ & new_n6746_;
  assign new_n6750_ = new_n6747_ | new_n6745_;
  assign new_n6751_ = new_n6749_ & new_n9743_;
  assign new_n6752_ = new_n6750_ | new_n9775_;
  assign new_n6753_ = new_n6752_ & new_n6743_;
  assign new_n6754_ = new_n6751_ | new_n6744_;
  assign new_n6755_ = new_n10150_ & new_n10151_;
  assign new_n6756_ = new_n10152_ | new_n10153_;
  assign new_n6757_ = new_n10152_ & new_n10153_;
  assign new_n6758_ = new_n10150_ | new_n10151_;
  assign new_n6759_ = new_n6758_ & new_n6756_;
  assign new_n6760_ = new_n6757_ | new_n6755_;
  assign new_n6761_ = new_n9548_ & new_n10154_;
  assign new_n6762_ = new_n9558_ | new_n10157_;
  assign new_n6763_ = new_n9570_ & new_n10157_;
  assign new_n6764_ = new_n9576_ | new_n10154_;
  assign new_n6765_ = new_n6764_ & new_n6762_;
  assign new_n6766_ = new_n6763_ | new_n6761_;
  assign new_n6767_ = new_n9581_ & new_n10159_;
  assign new_n6768_ = new_n9590_ | new_n10162_;
  assign new_n6769_ = new_n9598_ & new_n10162_;
  assign new_n6770_ = new_n9604_ | new_n10159_;
  assign new_n6771_ = new_n6770_ & new_n6768_;
  assign new_n6772_ = new_n6769_ | new_n6767_;
  assign new_n6773_ = new_n10164_ & new_n10165_;
  assign new_n6774_ = new_n10166_ | new_n10167_;
  assign new_n6775_ = new_n10166_ & new_n10167_;
  assign new_n6776_ = new_n10164_ | new_n10165_;
  assign new_n6777_ = new_n6776_ & new_n6774_;
  assign new_n6778_ = new_n6775_ | new_n6773_;
  assign new_n6779_ = new_n6778_ | new_n6759_;
  assign new_n6780_ = new_n6777_ | new_n6760_;
  assign new_n6781_ = new_n6780_ & new_n6779_;
  assign new_n6782_ = new_n10057_ & new_n9932_;
  assign new_n6783_ = new_n10062_ | new_n10036_;
  assign new_n6784_ = new_n6782_ & new_n9980_;
  assign new_n6785_ = new_n6783_ | new_n9985_;
  assign new_n6786_ = new_n10070_ & new_n9932_;
  assign new_n6787_ = new_n10075_ | new_n10037_;
  assign new_n6788_ = new_n6786_ & new_n9986_;
  assign new_n6789_ = new_n6787_ | new_n9979_;
  assign new_n6790_ = new_n6789_ & new_n6785_;
  assign new_n6791_ = new_n6788_ | new_n6784_;
  assign new_n6792_ = new_n10081_ & new_n9981_;
  assign new_n6793_ = new_n10090_ | new_n9986_;
  assign new_n6794_ = new_n10101_ & new_n9987_;
  assign new_n6795_ = new_n10109_ | new_n9981_;
  assign new_n6796_ = new_n6795_ & new_n6793_;
  assign new_n6797_ = new_n6794_ | new_n6792_;
  assign new_n6798_ = new_n6796_ & new_n10037_;
  assign new_n6799_ = new_n6797_ | new_n9933_;
  assign new_n6800_ = new_n6799_ & new_n6790_;
  assign new_n6801_ = new_n6798_ | new_n6791_;
  assign new_n6802_ = new_n10058_ & new_n9954_;
  assign new_n6803_ = new_n10064_ | new_n10043_;
  assign new_n6804_ = new_n6802_ & new_n4287_;
  assign new_n6805_ = new_n6803_ | new_n4286_;
  assign new_n6806_ = new_n10071_ & new_n9954_;
  assign new_n6807_ = new_n10077_ | new_n10044_;
  assign new_n6808_ = new_n6806_ & new_n4572_;
  assign new_n6809_ = new_n6807_ | new_n4573_;
  assign new_n6810_ = new_n6809_ & new_n6805_;
  assign new_n6811_ = new_n6808_ | new_n6804_;
  assign new_n6812_ = new_n10083_ & new_n10168_;
  assign new_n6813_ = new_n10090_ | new_n10169_;
  assign new_n6814_ = new_n10103_ & new_n10169_;
  assign new_n6815_ = new_n10109_ | new_n10168_;
  assign new_n6816_ = new_n6815_ & new_n6813_;
  assign new_n6817_ = new_n6814_ | new_n6812_;
  assign new_n6818_ = new_n6816_ & new_n10044_;
  assign new_n6819_ = new_n6817_ | new_n9955_;
  assign new_n6820_ = new_n6819_ & new_n6810_;
  assign new_n6821_ = new_n6818_ | new_n6811_;
  assign new_n6822_ = new_n10058_ & new_n9946_;
  assign new_n6823_ = new_n10064_ | new_n10040_;
  assign new_n6824_ = new_n6822_ & new_n4285_;
  assign new_n6825_ = new_n6823_ | new_n4284_;
  assign new_n6826_ = new_n10071_ & new_n9946_;
  assign new_n6827_ = new_n10077_ | new_n10041_;
  assign new_n6828_ = new_n6826_ & new_n4570_;
  assign new_n6829_ = new_n6827_ | new_n4571_;
  assign new_n6830_ = new_n6829_ & new_n6825_;
  assign new_n6831_ = new_n6828_ | new_n6824_;
  assign new_n6832_ = new_n10083_ & new_n10170_;
  assign new_n6833_ = new_n10092_ | new_n10171_;
  assign new_n6834_ = new_n10103_ & new_n10171_;
  assign new_n6835_ = new_n10111_ | new_n10170_;
  assign new_n6836_ = new_n6835_ & new_n6833_;
  assign new_n6837_ = new_n6834_ | new_n6832_;
  assign new_n6838_ = new_n6836_ & new_n10041_;
  assign new_n6839_ = new_n6837_ | new_n9947_;
  assign new_n6840_ = new_n6839_ & new_n6830_;
  assign new_n6841_ = new_n6838_ | new_n6831_;
  assign new_n6842_ = new_n10172_ & new_n10173_;
  assign new_n6843_ = new_n10174_ | new_n10175_;
  assign new_n6844_ = new_n10174_ & new_n10175_;
  assign new_n6845_ = new_n10172_ | new_n10173_;
  assign new_n6846_ = new_n6845_ & new_n6843_;
  assign new_n6847_ = new_n6844_ | new_n6842_;
  assign new_n6848_ = new_n4527_ & new_n4525_;
  assign new_n6849_ = new_n4526_ | new_n4524_;
  assign new_n6850_ = new_n10084_ & new_n4293_;
  assign new_n6851_ = new_n10092_ | new_n4292_;
  assign new_n6852_ = new_n4580_ & new_n10104_;
  assign new_n6853_ = new_n4581_ | new_n10111_;
  assign new_n6854_ = new_n6853_ & new_n6851_;
  assign new_n6855_ = new_n6852_ | new_n6850_;
  assign new_n6856_ = new_n6854_ & new_n10038_;
  assign new_n6857_ = new_n6855_ | new_n9939_;
  assign new_n6858_ = new_n6857_ & new_n6848_;
  assign new_n6859_ = new_n6856_ | new_n6849_;
  assign new_n6860_ = new_n4533_ & new_n4531_;
  assign new_n6861_ = new_n4532_ | new_n4530_;
  assign new_n6862_ = new_n10084_ & new_n4303_;
  assign new_n6863_ = new_n10093_ | new_n4302_;
  assign new_n6864_ = new_n4590_ & new_n10104_;
  assign new_n6865_ = new_n4591_ | new_n10112_;
  assign new_n6866_ = new_n6865_ & new_n6863_;
  assign new_n6867_ = new_n6864_ | new_n6862_;
  assign new_n6868_ = new_n6866_ & new_n9680_;
  assign new_n6869_ = new_n6867_ | new_n9677_;
  assign new_n6870_ = new_n6869_ & new_n6860_;
  assign new_n6871_ = new_n6868_ | new_n6861_;
  assign new_n6872_ = new_n10176_ & new_n10177_;
  assign new_n6873_ = new_n10178_ | new_n10179_;
  assign new_n6874_ = new_n10178_ & new_n10179_;
  assign new_n6875_ = new_n10176_ | new_n10177_;
  assign new_n6876_ = new_n6875_ & new_n6873_;
  assign new_n6877_ = new_n6874_ | new_n6872_;
  assign new_n6878_ = new_n10180_ | new_n10181_;
  assign new_n6879_ = new_n6878_ | new_n10182_;
  assign new_n6880_ = new_n10180_ | new_n10183_;
  assign new_n6881_ = new_n6880_ | new_n10184_;
  assign new_n6882_ = new_n6881_ & new_n6879_;
  assign new_n6883_ = new_n10185_ | new_n10183_;
  assign new_n6884_ = new_n6883_ | new_n10182_;
  assign new_n6885_ = new_n10185_ | new_n10181_;
  assign new_n6886_ = new_n6885_ | new_n10184_;
  assign new_n6887_ = new_n6886_ & new_n6884_;
  assign new_n6888_ = new_n6887_ & new_n6882_;
  assign new_n6889_ = new_n9548_ & new_n9974_;
  assign new_n6890_ = new_n9560_ | new_n10052_;
  assign new_n6891_ = new_n6889_ & new_n4291_;
  assign new_n6892_ = new_n6890_ | new_n4290_;
  assign new_n6893_ = new_n9570_ & new_n9974_;
  assign new_n6894_ = new_n9576_ | new_n10053_;
  assign new_n6895_ = new_n6893_ & new_n4576_;
  assign new_n6896_ = new_n6894_ | new_n4577_;
  assign new_n6897_ = new_n6896_ & new_n6892_;
  assign new_n6898_ = new_n6895_ | new_n6891_;
  assign new_n6899_ = new_n9583_ & new_n10186_;
  assign new_n6900_ = new_n9590_ | new_n10187_;
  assign new_n6901_ = new_n9600_ & new_n10187_;
  assign new_n6902_ = new_n9606_ | new_n10186_;
  assign new_n6903_ = new_n6902_ & new_n6900_;
  assign new_n6904_ = new_n6901_ | new_n6899_;
  assign new_n6905_ = new_n6903_ & new_n10053_;
  assign new_n6906_ = new_n6904_ | new_n9975_;
  assign new_n6907_ = new_n6906_ & new_n6897_;
  assign new_n6908_ = new_n6905_ | new_n6898_;
  assign new_n6909_ = new_n9549_ & new_n9967_;
  assign new_n6910_ = new_n9560_ | new_n10049_;
  assign new_n6911_ = new_n6909_ & new_n4289_;
  assign new_n6912_ = new_n6910_ | new_n4288_;
  assign new_n6913_ = new_n9569_ & new_n9967_;
  assign new_n6914_ = new_n9577_ | new_n10050_;
  assign new_n6915_ = new_n6913_ & new_n4574_;
  assign new_n6916_ = new_n6914_ | new_n4575_;
  assign new_n6917_ = new_n6916_ & new_n6912_;
  assign new_n6918_ = new_n6915_ | new_n6911_;
  assign new_n6919_ = new_n9583_ & new_n10188_;
  assign new_n6920_ = new_n9592_ | new_n10189_;
  assign new_n6921_ = new_n9600_ & new_n10189_;
  assign new_n6922_ = new_n9606_ | new_n10188_;
  assign new_n6923_ = new_n6922_ & new_n6920_;
  assign new_n6924_ = new_n6921_ | new_n6919_;
  assign new_n6925_ = new_n6923_ & new_n10050_;
  assign new_n6926_ = new_n6924_ | new_n9968_;
  assign new_n6927_ = new_n6926_ & new_n6917_;
  assign new_n6928_ = new_n6925_ | new_n6918_;
  assign new_n6929_ = new_n10190_ & new_n10191_;
  assign new_n6930_ = new_n10192_ | new_n10193_;
  assign new_n6931_ = new_n10192_ & new_n10193_;
  assign new_n6932_ = new_n10190_ | new_n10191_;
  assign new_n6933_ = new_n6932_ & new_n6930_;
  assign new_n6934_ = new_n6931_ | new_n6929_;
  assign new_n6935_ = new_n9549_ & new_n9959_;
  assign new_n6936_ = new_n9561_ | new_n10046_;
  assign new_n6937_ = new_n9592_ & new_n10045_;
  assign new_n6938_ = new_n9584_ | new_n9961_;
  assign new_n6939_ = new_n6938_ & new_n6936_;
  assign new_n6940_ = new_n6937_ | new_n6935_;
  assign new_n6941_ = new_n4537_ & new_n4535_;
  assign new_n6942_ = new_n4536_ | new_n4534_;
  assign new_n6943_ = new_n9584_ & new_n4305_;
  assign new_n6944_ = new_n9593_ | new_n4304_;
  assign new_n6945_ = new_n4592_ & new_n9599_;
  assign new_n6946_ = new_n4593_ | new_n9607_;
  assign new_n6947_ = new_n6946_ & new_n6944_;
  assign new_n6948_ = new_n6945_ | new_n6943_;
  assign new_n6949_ = new_n6947_ & new_n9690_;
  assign new_n6950_ = new_n6948_ | new_n9687_;
  assign new_n6951_ = new_n6950_ & new_n6941_;
  assign new_n6952_ = new_n6949_ | new_n6942_;
  assign new_n6953_ = new_n10194_ & new_n10195_;
  assign new_n6954_ = new_n10196_ | new_n10197_;
  assign new_n6955_ = new_n10196_ & new_n10197_;
  assign new_n6956_ = new_n10194_ | new_n10195_;
  assign new_n6957_ = new_n6956_ & new_n6954_;
  assign new_n6958_ = new_n6955_ | new_n6953_;
  assign new_n6959_ = new_n10198_ & new_n10199_;
  assign new_n6960_ = new_n6959_ & new_n10200_;
  assign new_n6961_ = new_n10198_ & new_n10202_;
  assign new_n6962_ = new_n6961_ & new_n10203_;
  assign new_n6963_ = new_n6962_ | new_n6960_;
  assign new_n6964_ = new_n10204_ & new_n10202_;
  assign new_n6965_ = new_n6964_ & new_n10200_;
  assign new_n6966_ = new_n10204_ & new_n10199_;
  assign new_n6967_ = new_n6966_ & new_n10203_;
  assign new_n6968_ = new_n6967_ | new_n6965_;
  assign new_n6969_ = new_n6968_ | new_n6963_;
  assign new_n6970_ = new_n10206_ & new_n10208_;
  assign new_n6971_ = new_n10210_ & new_n10212_;
  assign new_n6972_ = new_n4639_ & new_n4541_;
  assign new_n6973_ = new_n4638_ | new_n10213_;
  assign new_n6974_ = new_n6972_ & new_n4625_;
  assign new_n6975_ = new_n6973_ | new_n4624_;
  assign new_n6976_ = new_n6974_ & new_n4629_;
  assign new_n6977_ = new_n6975_ | new_n4628_;
  assign new_n6978_ = new_n6976_ & new_n4633_;
  assign new_n6979_ = new_n6977_ | new_n4632_;
  assign new_n6980_ = new_n4648_ & new_n4645_;
  assign new_n6981_ = new_n4649_ | new_n4644_;
  assign new_n6982_ = new_n10214_ & new_n10215_;
  assign new_n6983_ = new_n10216_ | new_n10217_;
  assign new_n6984_ = new_n10216_ & new_n10217_;
  assign new_n6985_ = new_n10214_ | new_n10215_;
  assign new_n6986_ = new_n6985_ & new_n6983_;
  assign new_n6987_ = new_n6984_ | new_n6982_;
  assign new_n6988_ = new_n10218_ & new_n10220_;
  assign new_n6989_ = new_n10222_ | new_n10225_;
  assign new_n6990_ = new_n10222_ & new_n10225_;
  assign new_n6991_ = new_n10218_ | new_n10220_;
  assign new_n6992_ = new_n6991_ & new_n6989_;
  assign new_n6993_ = new_n6990_ | new_n6988_;
  assign new_n6994_ = new_n6993_ | new_n10228_;
  assign new_n6995_ = new_n6992_ | new_n10229_;
  assign new_n6996_ = new_n6995_ & new_n6994_;
  assign new_n6997_ = new_n4641_ & new_n4539_;
  assign new_n6998_ = new_n4640_ | new_n10230_;
  assign new_n6999_ = new_n6997_ & new_n4627_;
  assign new_n7000_ = new_n6998_ | new_n4626_;
  assign new_n7001_ = new_n6999_ & new_n4635_;
  assign new_n7002_ = new_n7000_ | new_n4634_;
  assign new_n7003_ = new_n7001_ & new_n4637_;
  assign new_n7004_ = new_n7002_ | new_n4636_;
  assign new_n7005_ = new_n4647_ & new_n4643_;
  assign new_n7006_ = new_n4646_ | new_n4642_;
  assign new_n7007_ = new_n10231_ & new_n10232_;
  assign new_n7008_ = new_n10233_ | new_n10234_;
  assign new_n7009_ = new_n10233_ & new_n10234_;
  assign new_n7010_ = new_n10231_ | new_n10232_;
  assign new_n7011_ = new_n7010_ & new_n7008_;
  assign new_n7012_ = new_n7009_ | new_n7007_;
  assign new_n7013_ = new_n10235_ & new_n10238_;
  assign new_n7014_ = new_n10240_ | new_n10242_;
  assign new_n7015_ = new_n10240_ & new_n10242_;
  assign new_n7016_ = new_n10235_ | new_n10238_;
  assign new_n7017_ = new_n7016_ & new_n7014_;
  assign new_n7018_ = new_n7015_ | new_n7013_;
  assign new_n7019_ = new_n7018_ | new_n10245_;
  assign new_n7020_ = new_n7017_ | new_n10246_;
  assign new_n7021_ = new_n7020_ & new_n7019_;
  assign new_n7022_ = new_n10248_ & new_n10250_;
  assign new_n7023_ = new_n10252_ | new_n4543_;
  assign new_n7024_ = new_n10255_ & new_n10260_;
  assign new_n7025_ = new_n10262_ | new_n10264_;
  assign new_n7026_ = new_n7024_ & new_n10248_;
  assign new_n7027_ = new_n7025_ | new_n10252_;
  assign new_n7028_ = new_n10266_ & new_n10255_;
  assign new_n7029_ = new_n10269_ | new_n10262_;
  assign new_n7030_ = new_n7028_ & new_n10249_;
  assign new_n7031_ = new_n7029_ | new_n10251_;
  assign new_n7032_ = new_n7023_ & new_n6282_;
  assign new_n7033_ = new_n7022_ | new_n10270_;
  assign new_n7034_ = new_n7032_ & new_n7027_;
  assign new_n7035_ = new_n7033_ | new_n7026_;
  assign new_n7036_ = new_n10272_ & new_n7031_;
  assign new_n7037_ = new_n10274_ | new_n7030_;
  assign new_n7038_ = new_n10276_ & new_n4651_;
  assign new_n7039_ = new_n10278_ | new_n4650_;
  assign new_n7040_ = new_n4241_ & new_n4235_;
  assign new_n7041_ = new_n10279_ | new_n10280_;
  assign new_n7042_ = new_n10281_ & new_n10282_;
  assign new_n7043_ = new_n10283_ | new_n10284_;
  assign new_n7044_ = new_n10283_ & new_n10284_;
  assign new_n7045_ = new_n10281_ | new_n10282_;
  assign new_n7046_ = new_n7045_ & new_n7043_;
  assign new_n7047_ = new_n7044_ | new_n7042_;
  assign new_n7048_ = new_n10285_ & new_n10286_;
  assign new_n7049_ = new_n10287_ | new_n10288_;
  assign new_n7050_ = new_n10287_ & new_n10288_;
  assign new_n7051_ = new_n10285_ | new_n10286_;
  assign new_n7052_ = new_n7051_ & new_n7049_;
  assign new_n7053_ = new_n7050_ | new_n7048_;
  assign new_n7054_ = new_n7052_ & new_n10269_;
  assign new_n7055_ = new_n7053_ & new_n10266_;
  assign new_n7056_ = new_n7055_ | new_n7054_;
  assign new_n7057_ = new_n10276_ & new_n10260_;
  assign new_n7058_ = new_n10278_ | new_n10264_;
  assign new_n7059_ = new_n10277_ & new_n10263_;
  assign new_n7060_ = new_n10275_ | new_n10261_;
  assign new_n7061_ = new_n7060_ & new_n7058_;
  assign new_n7062_ = new_n7059_ | new_n7057_;
  assign new_n7063_ = new_n10289_ & new_n10272_;
  assign new_n7064_ = new_n10290_ | new_n10274_;
  assign new_n7065_ = new_n10290_ & new_n10273_;
  assign new_n7066_ = new_n10289_ | new_n10271_;
  assign new_n7067_ = new_n7066_ & new_n7064_;
  assign new_n7068_ = new_n7065_ | new_n7063_;
  assign new_n7069_ = new_n7067_ & new_n10268_;
  assign new_n7070_ = new_n7068_ & new_n10267_;
  assign new_n7071_ = new_n7070_ | new_n7069_;
  assign new_n7072_ = new_n10292_ & new_n10294_;
  assign new_n7073_ = new_n10297_ | new_n4545_;
  assign new_n7074_ = new_n10303_ & new_n10308_;
  assign new_n7075_ = new_n10310_ | new_n10312_;
  assign new_n7076_ = new_n7074_ & new_n10292_;
  assign new_n7077_ = new_n7075_ | new_n10297_;
  assign new_n7078_ = new_n10314_ & new_n10303_;
  assign new_n7079_ = new_n10317_ | new_n10310_;
  assign new_n7080_ = new_n7078_ & new_n10293_;
  assign new_n7081_ = new_n7079_ | new_n10298_;
  assign new_n7082_ = new_n7073_ & new_n10298_;
  assign new_n7083_ = new_n7072_ | new_n10293_;
  assign new_n7084_ = new_n7082_ & new_n7077_;
  assign new_n7085_ = new_n7083_ | new_n7076_;
  assign new_n7086_ = new_n10319_ & new_n7081_;
  assign new_n7087_ = new_n10321_ | new_n7080_;
  assign new_n7088_ = new_n10323_ & new_n4653_;
  assign new_n7089_ = new_n10325_ | new_n4652_;
  assign new_n7090_ = new_n4239_ & new_n4237_;
  assign new_n7091_ = new_n10326_ | new_n10327_;
  assign new_n7092_ = new_n10328_ & new_n10329_;
  assign new_n7093_ = new_n10330_ | new_n10331_;
  assign new_n7094_ = new_n10330_ & new_n10331_;
  assign new_n7095_ = new_n10328_ | new_n10329_;
  assign new_n7096_ = new_n7095_ & new_n7093_;
  assign new_n7097_ = new_n7094_ | new_n7092_;
  assign new_n7098_ = new_n10332_ & new_n10333_;
  assign new_n7099_ = new_n10334_ | new_n10335_;
  assign new_n7100_ = new_n10334_ & new_n10335_;
  assign new_n7101_ = new_n10332_ | new_n10333_;
  assign new_n7102_ = new_n7101_ & new_n7099_;
  assign new_n7103_ = new_n7100_ | new_n7098_;
  assign new_n7104_ = new_n7103_ | new_n10314_;
  assign new_n7105_ = new_n7102_ | new_n10317_;
  assign new_n7106_ = new_n7105_ & new_n7104_;
  assign new_n7107_ = new_n10323_ & new_n10308_;
  assign new_n7108_ = new_n10325_ | new_n10312_;
  assign new_n7109_ = new_n10324_ & new_n10311_;
  assign new_n7110_ = new_n10322_ | new_n10309_;
  assign new_n7111_ = new_n7110_ & new_n7108_;
  assign new_n7112_ = new_n7109_ | new_n7107_;
  assign new_n7113_ = new_n10336_ & new_n10319_;
  assign new_n7114_ = new_n10337_ | new_n10321_;
  assign new_n7115_ = new_n10337_ & new_n10320_;
  assign new_n7116_ = new_n10336_ | new_n10318_;
  assign new_n7117_ = new_n7116_ & new_n7114_;
  assign new_n7118_ = new_n7115_ | new_n7113_;
  assign new_n7119_ = new_n7118_ | new_n10315_;
  assign new_n7120_ = new_n7117_ | new_n10316_;
  assign new_n7121_ = new_n7120_ & new_n7119_;
  assign new_n7122_ = new_n9830_ & new_n10338_;
  assign new_n7123_ = new_n9835_ & new_n3392_;
  assign new_n7124_ = new_n7123_ | new_n7122_;
  assign new_n7125_ = new_n10340_ & new_n10342_;
  assign new_n7126_ = new_n10344_ | new_n10346_;
  assign new_n7127_ = new_n10344_ & new_n10346_;
  assign new_n7128_ = new_n10340_ | new_n10342_;
  assign new_n7129_ = new_n7128_ & new_n7126_;
  assign new_n7130_ = new_n7127_ | new_n7125_;
  assign new_n7131_ = new_n6365_ & new_n10348_;
  assign new_n7132_ = new_n10350_ & new_n3551_;
  assign new_n7133_ = new_n7132_ | new_n7131_;
  assign new_n7134_ = new_n6377_ & new_n10352_;
  assign new_n7135_ = new_n10354_ & new_n3579_;
  assign new_n7136_ = new_n7135_ | new_n7134_;
  assign new_n7137_ = new_n6371_ & new_n10356_;
  assign new_n7138_ = new_n10358_ & new_n3583_;
  assign new_n7139_ = new_n7138_ | new_n7137_;
  assign new_n7140_ = new_n10360_ & new_n10362_;
  assign new_n7141_ = new_n7140_ & new_n4129_;
  assign new_n7142_ = new_n10360_ & new_n10364_;
  assign new_n7143_ = new_n7142_ & new_n10366_;
  assign new_n7144_ = new_n9917_ & new_n10362_;
  assign new_n7145_ = new_n7144_ & new_n9711_;
  assign new_n7146_ = new_n9918_ & new_n10364_;
  assign new_n7147_ = new_n7146_ & new_n9709_;
  assign new_n7148_ = new_n9921_ & new_n10361_;
  assign new_n7149_ = new_n7148_ & new_n9704_;
  assign new_n7150_ = new_n9922_ & new_n10363_;
  assign new_n7151_ = new_n7150_ & new_n9702_;
  assign new_n7152_ = new_n10339_ | new_n10345_;
  assign new_n7153_ = new_n10350_ & new_n10348_;
  assign new_n7154_ = new_n10354_ & new_n10352_;
  assign new_n7155_ = new_n10358_ & new_n10356_;
  assign new_n7156_ = new_n10369_ & new_n10370_;
  assign new_n7157_ = new_n10371_ & new_n10372_;
  assign new_n7158_ = new_n10373_ | new_n10374_;
  assign new_n7159_ = new_n10373_ & new_n10374_;
  assign new_n7160_ = new_n10371_ | new_n10372_;
  assign new_n7161_ = new_n7160_ & new_n7158_;
  assign new_n7162_ = new_n7159_ | new_n7157_;
  assign new_n7163_ = new_n10375_ & new_n10221_;
  assign new_n7164_ = new_n10376_ | new_n10224_;
  assign new_n7165_ = new_n10376_ & new_n10226_;
  assign new_n7166_ = new_n10375_ | new_n10221_;
  assign new_n7167_ = new_n7166_ & new_n7164_;
  assign new_n7168_ = new_n7165_ | new_n7163_;
  assign new_n7169_ = new_n7167_ & new_n10229_;
  assign new_n7170_ = new_n7168_ & new_n10228_;
  assign new_n7171_ = new_n7170_ | new_n7169_;
  assign new_n7172_ = new_n10377_ & new_n10380_;
  assign new_n7173_ = new_n10382_ & new_n10383_;
  assign new_n7174_ = new_n10384_ | new_n10385_;
  assign new_n7175_ = new_n10384_ & new_n10385_;
  assign new_n7176_ = new_n10382_ | new_n10383_;
  assign new_n7177_ = new_n7176_ & new_n7174_;
  assign new_n7178_ = new_n7175_ | new_n7173_;
  assign new_n7179_ = new_n10386_ & new_n10237_;
  assign new_n7180_ = new_n10387_ | new_n10243_;
  assign new_n7181_ = new_n10387_ & new_n10243_;
  assign new_n7182_ = new_n10386_ | new_n10239_;
  assign new_n7183_ = new_n7182_ & new_n7180_;
  assign new_n7184_ = new_n7181_ | new_n7179_;
  assign new_n7185_ = new_n7183_ & new_n10246_;
  assign new_n7186_ = new_n7184_ & new_n10245_;
  assign new_n7187_ = new_n7186_ | new_n7185_;
  assign new_n7188_ = new_n10388_ & new_n10391_;
  assign new_n7189_ = new_n10369_ | new_n10370_;
  assign new_n7190_ = new_n10377_ | new_n10380_;
  assign new_n7191_ = new_n10388_ | new_n10391_;
  assign new_n7192_ = new_n9699_ & new_n10393_;
  assign new_n7193_ = new_n9705_ & new_n10394_;
  assign new_n7194_ = new_n7193_ | new_n7192_;
  assign new_n7195_ = new_n6552_ & new_n10208_;
  assign new_n7196_ = new_n10206_ & new_n3559_;
  assign new_n7197_ = new_n7196_ | new_n7195_;
  assign new_n7198_ = new_n6546_ & new_n10212_;
  assign new_n7199_ = new_n10210_ & new_n3587_;
  assign new_n7200_ = new_n7199_ | new_n7198_;
  assign new_n7201_ = new_n9824_ & new_n3480_;
  assign new_n7202_ = new_n10396_ & new_n10399_;
  assign new_n7203_ = new_n10401_ | new_n10402_;
  assign new_n7204_ = new_n10403_ & new_n10406_;
  assign new_n7205_ = new_n10409_ & new_n10411_;
  assign new_n7206_ = new_n10413_ | new_n10414_;
  assign new_n7207_ = new_n10415_ | new_n10417_;
  assign new_n7208_ = new_n10421_ & new_n10396_;
  assign new_n7209_ = new_n10425_ | new_n10401_;
  assign new_n7210_ = new_n7208_ & new_n10428_;
  assign new_n7211_ = new_n7209_ | new_n10431_;
  assign new_n7212_ = new_n10433_ & new_n10406_;
  assign new_n7213_ = new_n9819_ & new_n10434_;
  assign new_n7214_ = new_n10436_ & new_n10397_;
  assign new_n7215_ = new_n6355_ | new_n10400_;
  assign new_n7216_ = new_n10437_ & new_n10405_;
  assign new_n7217_ = new_n7216_ & new_n10421_;
  assign new_n7218_ = new_n10439_ & new_n10409_;
  assign new_n7219_ = new_n10441_ | new_n10413_;
  assign new_n7220_ = new_n7218_ & new_n10444_;
  assign new_n7221_ = new_n7219_ | new_n10448_;
  assign new_n7222_ = new_n10453_ | new_n10417_;
  assign new_n7223_ = new_n10412_ | new_n10448_;
  assign new_n7224_ = new_n10454_ | new_n10418_;
  assign new_n7225_ = new_n7224_ | new_n10441_;
  assign new_n7226_ = new_n10407_ & new_n10456_;
  assign new_n7227_ = new_n10418_ | new_n10457_;
  assign new_n7228_ = new_n10454_ | new_n10442_;
  assign new_n7229_ = new_n10415_ & new_n10457_;
  assign new_n7230_ = new_n7205_ | new_n10458_;
  assign new_n7231_ = new_n7229_ & new_n10453_;
  assign new_n7232_ = new_n7230_ | new_n7220_;
  assign new_n7233_ = new_n10460_ & new_n7228_;
  assign new_n7234_ = new_n10439_ & new_n10444_;
  assign new_n7235_ = new_n10442_ | new_n10449_;
  assign new_n7236_ = new_n7235_ & new_n10414_;
  assign new_n7237_ = new_n10461_ | new_n10411_;
  assign new_n7238_ = new_n10462_ | new_n10461_;
  assign new_n7239_ = new_n10463_ | new_n10464_;
  assign new_n7240_ = new_n10422_ & new_n10428_;
  assign new_n7241_ = new_n10425_ | new_n10431_;
  assign new_n7242_ = new_n7241_ & new_n10402_;
  assign new_n7243_ = new_n7240_ | new_n10399_;
  assign new_n7244_ = new_n10436_ & new_n10422_;
  assign new_n7245_ = new_n7244_ | new_n10465_;
  assign new_n7246_ = new_n10437_ & new_n10423_;
  assign new_n7247_ = new_n7215_ | new_n10424_;
  assign new_n7248_ = new_n7203_ & new_n6348_;
  assign new_n7249_ = new_n10403_ | new_n10456_;
  assign new_n7250_ = new_n7248_ & new_n7211_;
  assign new_n7251_ = new_n7249_ | new_n10433_;
  assign new_n7252_ = new_n10467_ & new_n7247_;
  assign new_n7253_ = new_n10469_ | new_n7246_;
  assign new_n7254_ = new_n9786_ & new_n9789_;
  assign new_n7255_ = new_n9779_ | new_n9783_;
  assign new_n7256_ = new_n7254_ | new_n7252_;
  assign new_n7257_ = new_n7255_ | new_n7253_;
  assign new_n7258_ = new_n7257_ & new_n7256_;
  assign new_n7259_ = new_n10470_ & new_n10471_;
  assign new_n7260_ = new_n10463_ & new_n10464_;
  assign new_n7261_ = new_n10470_ | new_n10471_;
  assign new_n7262_ = new_n10472_ & new_n10474_;
  assign new_n7263_ = new_n10475_ & new_n10477_;
  assign new_n7264_ = new_n10478_ | new_n10479_;
  assign new_n7265_ = new_n7264_ | new_n10480_;
  assign new_n7266_ = new_n7265_ | new_n10481_;
  assign new_n7267_ = new_n10482_ & new_n10483_;
  assign new_n7268_ = new_n7267_ & new_n10484_;
  assign new_n7269_ = new_n7268_ & new_n10485_;
  assign new_n7270_ = new_n10474_ & new_n10486_;
  assign new_n7271_ = new_n7270_ | new_n10487_;
  assign new_n7272_ = new_n10477_ & new_n10488_;
  assign new_n7273_ = new_n7272_ | new_n10489_;
  assign new_n7274_ = new_n10467_ & new_n10427_;
  assign new_n7275_ = new_n10469_ | new_n10432_;
  assign new_n7276_ = new_n10468_ & new_n10432_;
  assign new_n7277_ = new_n10466_ | new_n10429_;
  assign new_n7278_ = new_n7277_ & new_n7275_;
  assign new_n7279_ = new_n7276_ | new_n7274_;
  assign new_n7280_ = new_n7279_ | new_n10465_;
  assign new_n7281_ = new_n7278_ | new_n7242_;
  assign new_n7282_ = new_n7281_ & new_n7280_;
  assign new_n7283_ = new_n10460_ & new_n10445_;
  assign new_n7284_ = new_n10490_ | new_n10449_;
  assign new_n7285_ = new_n10490_ & new_n10451_;
  assign new_n7286_ = new_n10459_ | new_n10445_;
  assign new_n7287_ = new_n7286_ & new_n7284_;
  assign new_n7288_ = new_n7285_ | new_n7283_;
  assign new_n7289_ = new_n7287_ & new_n7236_;
  assign new_n7290_ = new_n7288_ & new_n10462_;
  assign new_n7291_ = new_n7290_ | new_n7289_;
  assign new_n7292_ = new_n10491_ & new_n10494_;
  assign new_n7293_ = new_n10496_ & new_n10497_;
  assign new_n7294_ = new_n7293_ | new_n7292_;
  assign new_n7295_ = new_n10498_ & new_n10494_;
  assign new_n7296_ = new_n10499_ & new_n10497_;
  assign new_n7297_ = new_n7296_ | new_n7295_;
  assign new_n7298_ = new_n10502_ & new_n10505_;
  assign new_n7299_ = new_n10507_ & new_n2538_;
  assign new_n7300_ = new_n7299_ | new_n7298_;
  assign new_n7301_ = new_n10502_ & new_n10508_;
  assign new_n7302_ = new_n10507_ & new_n2542_;
  assign new_n7303_ = new_n7302_ | new_n7301_;
  assign new_n7304_ = new_n10503_ & new_n10509_;
  assign new_n7305_ = new_n10506_ & new_n2546_;
  assign new_n7306_ = new_n7305_ | new_n7304_;
  assign G5193 = new_n8486_;
  assign G5194 = new_n8501_;
  assign G5195 = new_n8445_;
  assign G5196 = new_n10511_;
  assign G5197 = new_n3511_;
  assign G5198 = new_n3519_;
  assign G5199 = new_n4710_;
  assign G5200 = new_n3619_;
  assign G5201 = G5196;
  assign G5202 = new_n10510_;
  assign G5203 = new_n3507_;
  assign G5204 = new_n3515_;
  assign G5205 = new_n4711_;
  assign G5206 = new_n9477_;
  assign G5207 = new_n9471_;
  assign G5208 = new_n9473_;
  assign G5209 = new_n9470_;
  assign G5210 = new_n4712_;
  assign G5211 = new_n4713_;
  assign G5212 = new_n4714_;
  assign G5213 = new_n4715_;
  assign G5214 = new_n9331_;
  assign G5215 = new_n8443_;
  assign G5216 = new_n8444_;
  assign G5217 = new_n10512_;
  assign G5218 = new_n3474_;
  assign G5219 = G5217;
  assign G5220 = new_n4718_;
  assign G5221 = new_n8460_;
  assign G5222 = new_n10514_;
  assign G5223 = G5222;
  assign G5224 = new_n10515_;
  assign G5225 = G5224;
  assign G5226 = new_n10516_;
  assign G5227 = G5226;
  assign G5228 = new_n4722_;
  assign G5229 = new_n10517_;
  assign G5230 = G5229;
  assign G5231 = new_n4730_;
  assign G5232 = ~new_n4740_;
  assign G5233 = ~new_n4748_;
  assign G5234 = ~new_n4756_;
  assign G5235 = ~new_n4764_;
  assign G5236 = ~new_n4834_;
  assign G5237 = ~new_n4922_;
  assign G5238 = ~new_n4926_;
  assign G5239 = ~new_n4938_;
  assign G5240 = ~new_n4942_;
  assign G5241 = ~new_n4954_;
  assign G5242 = ~new_n9475_;
  assign G5243 = ~new_n9476_;
  assign G5244 = ~new_n5060_;
  assign G5245 = ~new_n5101_;
  assign G5246 = ~new_n5142_;
  assign G5247 = ~new_n5153_;
  assign G5248 = ~new_n8992_;
  assign G5249 = ~new_n9441_;
  assign G5250 = ~new_n9034_;
  assign G5251 = new_n9468_;
  assign G5252 = new_n5232_;
  assign G5253 = ~new_n9411_;
  assign G5254 = ~new_n9421_;
  assign G5255 = ~new_n9431_;
  assign G5256 = new_n5314_;
  assign G5257 = ~new_n9415_;
  assign G5258 = ~new_n9425_;
  assign G5259 = ~new_n9435_;
  assign G5260 = ~new_n9445_;
  assign G5261 = ~new_n9472_;
  assign G5262 = ~new_n9474_;
  assign G5263 = ~new_n5546_;
  assign G5264 = ~new_n5579_;
  assign G5265 = new_n5591_;
  assign G5266 = new_n5603_;
  assign G5267 = new_n5614_;
  assign G5268 = new_n5625_;
  assign G5269 = new_n5636_;
  assign G5270 = new_n5647_;
  assign G5271 = new_n5658_;
  assign G5272 = new_n5669_;
  assign G5273 = new_n5680_;
  assign G5274 = new_n5691_;
  assign G5275 = new_n5703_;
  assign G5276 = new_n5715_;
  assign G5277 = new_n5727_;
  assign G5278 = new_n5739_;
  assign G5279 = new_n5751_;
  assign G5280 = new_n5763_;
  assign G5281 = new_n5775_;
  assign G5282 = new_n5787_;
  assign G5283 = new_n5808_;
  assign G5284 = new_n5812_;
  assign G5285 = ~new_n9483_;
  assign G5286 = ~new_n9493_;
  assign G5287 = ~new_n9503_;
  assign G5288 = ~new_n9513_;
  assign G5289 = ~new_n5853_;
  assign G5290 = ~new_n9487_;
  assign G5291 = ~new_n9497_;
  assign G5292 = ~new_n9507_;
  assign G5293 = ~new_n9517_;
  assign G5294 = new_n5906_;
  assign G5295 = new_n5917_;
  assign G5296 = new_n5928_;
  assign G5297 = new_n5939_;
  assign G5298 = new_n5950_;
  assign G5299 = new_n5961_;
  assign G5300 = new_n5972_;
  assign G5301 = new_n5983_;
  assign G5302 = new_n5995_;
  assign G5303 = new_n6007_;
  assign G5304 = new_n6019_;
  assign G5305 = new_n6031_;
  assign G5306 = new_n6043_;
  assign G5307 = new_n6055_;
  assign G5308 = new_n6067_;
  assign G5309 = new_n6079_;
  assign G5310 = ~new_n6095_;
  assign G5311 = ~new_n6110_;
  assign G5312 = new_n6133_;
  assign G5313 = new_n6144_;
  assign G5314 = ~new_n6156_;
  assign G5315 = ~new_n6168_;
  assign n2610_li = new_n2328_;
  assign n2613_li = new_n2684_;
  assign n2616_li = new_n2686_;
  assign n2619_li = new_n2688_;
  assign n2622_li = new_n2330_;
  assign n2625_li = new_n2692_;
  assign n2628_li = new_n2694_;
  assign n2631_li = new_n2696_;
  assign n2634_li = new_n2332_;
  assign n2637_li = new_n2700_;
  assign n2640_li = new_n2702_;
  assign n2643_li = new_n2704_;
  assign n2646_li = new_n2334_;
  assign n2649_li = new_n2708_;
  assign n2652_li = new_n2710_;
  assign n2655_li = new_n2712_;
  assign n2658_li = new_n2336_;
  assign n2661_li = new_n2716_;
  assign n2664_li = new_n2718_;
  assign n2667_li = new_n2720_;
  assign n2670_li = new_n2338_;
  assign n2673_li = new_n2724_;
  assign n2676_li = new_n2726_;
  assign n2679_li = new_n2728_;
  assign n2682_li = new_n2340_;
  assign n2685_li = new_n2732_;
  assign n2688_li = new_n2734_;
  assign n2691_li = new_n2736_;
  assign n2694_li = new_n2342_;
  assign n2697_li = new_n2740_;
  assign n2700_li = new_n2742_;
  assign n2703_li = new_n2744_;
  assign n2706_li = new_n2344_;
  assign n2709_li = new_n2748_;
  assign n2712_li = new_n2750_;
  assign n2715_li = new_n2752_;
  assign n2718_li = new_n2346_;
  assign n2721_li = new_n2756_;
  assign n2724_li = new_n2758_;
  assign n2727_li = new_n2760_;
  assign n2730_li = new_n2348_;
  assign n2733_li = new_n2764_;
  assign n2736_li = new_n2766_;
  assign n2739_li = new_n2768_;
  assign n2742_li = new_n2350_;
  assign n2745_li = new_n2772_;
  assign n2748_li = new_n2774_;
  assign n2751_li = new_n2776_;
  assign n2754_li = new_n2352_;
  assign n2757_li = new_n2780_;
  assign n2760_li = new_n2782_;
  assign n2763_li = new_n2784_;
  assign n2766_li = new_n2354_;
  assign n2769_li = new_n2788_;
  assign n2772_li = new_n2790_;
  assign n2775_li = new_n2792_;
  assign n2778_li = new_n2356_;
  assign n2781_li = new_n2796_;
  assign n2784_li = new_n2798_;
  assign n2787_li = new_n2800_;
  assign n2790_li = new_n2358_;
  assign n2793_li = new_n2804_;
  assign n2796_li = new_n2806_;
  assign n2799_li = new_n2808_;
  assign n2802_li = new_n2360_;
  assign n2805_li = new_n2812_;
  assign n2808_li = new_n2814_;
  assign n2811_li = new_n2816_;
  assign n2814_li = new_n2362_;
  assign n2817_li = new_n2820_;
  assign n2820_li = new_n2822_;
  assign n2823_li = new_n2824_;
  assign n2826_li = new_n2364_;
  assign n2829_li = new_n2828_;
  assign n2832_li = new_n2830_;
  assign n2835_li = new_n2832_;
  assign n2838_li = new_n2366_;
  assign n2841_li = new_n2836_;
  assign n2844_li = new_n2838_;
  assign n2847_li = new_n2840_;
  assign n2850_li = new_n2368_;
  assign n2853_li = new_n2844_;
  assign n2856_li = new_n2846_;
  assign n2859_li = new_n2848_;
  assign n2862_li = new_n2370_;
  assign n2865_li = new_n2852_;
  assign n2868_li = new_n2854_;
  assign n2871_li = new_n2856_;
  assign n2874_li = new_n2372_;
  assign n2877_li = new_n2860_;
  assign n2880_li = new_n2862_;
  assign n2883_li = new_n2864_;
  assign n2886_li = new_n2374_;
  assign n2889_li = new_n2868_;
  assign n2892_li = new_n2870_;
  assign n2895_li = new_n2872_;
  assign n2898_li = new_n2376_;
  assign n2901_li = new_n2876_;
  assign n2904_li = new_n2878_;
  assign n2907_li = new_n2880_;
  assign n2910_li = new_n2378_;
  assign n2913_li = new_n2884_;
  assign n2916_li = new_n2886_;
  assign n2919_li = new_n2888_;
  assign n2922_li = new_n2380_;
  assign n2925_li = new_n2892_;
  assign n2928_li = new_n2894_;
  assign n2931_li = new_n2896_;
  assign n2934_li = new_n2382_;
  assign n2937_li = new_n2900_;
  assign n2940_li = new_n2902_;
  assign n2943_li = new_n2904_;
  assign n2946_li = new_n2384_;
  assign n2949_li = new_n2908_;
  assign n2952_li = new_n2910_;
  assign n2955_li = new_n2912_;
  assign n2958_li = new_n2386_;
  assign n2961_li = new_n2916_;
  assign n2964_li = new_n2918_;
  assign n2967_li = new_n2920_;
  assign n2970_li = new_n2388_;
  assign n2973_li = new_n2924_;
  assign n2976_li = new_n2926_;
  assign n2979_li = new_n2928_;
  assign n2982_li = new_n2390_;
  assign n2985_li = new_n2932_;
  assign n2988_li = new_n2934_;
  assign n2991_li = new_n2936_;
  assign n2994_li = new_n2392_;
  assign n2997_li = new_n2940_;
  assign n3000_li = new_n2942_;
  assign n3003_li = new_n2944_;
  assign n3006_li = new_n2394_;
  assign n3009_li = new_n2948_;
  assign n3012_li = new_n2950_;
  assign n3015_li = new_n2952_;
  assign n3018_li = new_n2396_;
  assign n3021_li = new_n2956_;
  assign n3024_li = new_n2958_;
  assign n3027_li = new_n2960_;
  assign n3030_li = new_n2398_;
  assign n3033_li = new_n2964_;
  assign n3036_li = new_n2966_;
  assign n3039_li = new_n2968_;
  assign n3042_li = new_n2400_;
  assign n3045_li = new_n2972_;
  assign n3048_li = new_n2974_;
  assign n3051_li = new_n2976_;
  assign n3054_li = new_n2402_;
  assign n3057_li = new_n2980_;
  assign n3060_li = new_n2982_;
  assign n3063_li = new_n2984_;
  assign n3066_li = new_n2404_;
  assign n3069_li = new_n2988_;
  assign n3072_li = new_n2990_;
  assign n3075_li = new_n2992_;
  assign n3078_li = new_n2406_;
  assign n3081_li = new_n2996_;
  assign n3084_li = new_n2998_;
  assign n3087_li = new_n3000_;
  assign n3090_li = new_n2408_;
  assign n3093_li = new_n3004_;
  assign n3096_li = new_n3006_;
  assign n3099_li = new_n3008_;
  assign n3102_li = new_n2410_;
  assign n3105_li = new_n3012_;
  assign n3108_li = new_n3014_;
  assign n3111_li = new_n3016_;
  assign n3114_li = new_n2412_;
  assign n3117_li = new_n3020_;
  assign n3120_li = new_n3022_;
  assign n3123_li = new_n3024_;
  assign n3126_li = new_n2414_;
  assign n3129_li = new_n3028_;
  assign n3132_li = new_n3030_;
  assign n3135_li = new_n3032_;
  assign n3138_li = new_n2416_;
  assign n3141_li = new_n3036_;
  assign n3144_li = new_n3038_;
  assign n3147_li = new_n3040_;
  assign n3150_li = new_n2418_;
  assign n3153_li = new_n3044_;
  assign n3156_li = new_n3046_;
  assign n3159_li = new_n3048_;
  assign n3162_li = new_n2420_;
  assign n3165_li = new_n3052_;
  assign n3168_li = new_n3054_;
  assign n3171_li = new_n3056_;
  assign n3174_li = new_n2422_;
  assign n3177_li = new_n3060_;
  assign n3180_li = new_n3062_;
  assign n3183_li = new_n3064_;
  assign n3186_li = new_n2424_;
  assign n3189_li = new_n3068_;
  assign n3192_li = new_n3070_;
  assign n3195_li = new_n3072_;
  assign n3198_li = new_n2426_;
  assign n3201_li = new_n3076_;
  assign n3204_li = new_n3078_;
  assign n3207_li = new_n3080_;
  assign n3210_li = new_n2428_;
  assign n3213_li = new_n3084_;
  assign n3216_li = new_n3086_;
  assign n3219_li = new_n3088_;
  assign n3222_li = new_n2430_;
  assign n3225_li = new_n3092_;
  assign n3228_li = new_n3094_;
  assign n3231_li = new_n3096_;
  assign n3234_li = new_n2432_;
  assign n3237_li = new_n3100_;
  assign n3240_li = new_n3102_;
  assign n3243_li = new_n3104_;
  assign n3246_li = new_n2434_;
  assign n3249_li = new_n3108_;
  assign n3252_li = new_n3110_;
  assign n3255_li = new_n3112_;
  assign n3258_li = new_n2436_;
  assign n3261_li = new_n3116_;
  assign n3264_li = new_n3118_;
  assign n3267_li = new_n3120_;
  assign n3270_li = new_n2438_;
  assign n3273_li = new_n3124_;
  assign n3276_li = new_n3126_;
  assign n3279_li = new_n3128_;
  assign n3282_li = new_n2440_;
  assign n3285_li = new_n3132_;
  assign n3288_li = new_n3134_;
  assign n3291_li = new_n3136_;
  assign n3294_li = new_n2442_;
  assign n3297_li = new_n3140_;
  assign n3300_li = new_n3142_;
  assign n3303_li = new_n3144_;
  assign n3306_li = new_n2444_;
  assign n3309_li = new_n3148_;
  assign n3312_li = new_n3150_;
  assign n3315_li = new_n3152_;
  assign n3318_li = new_n2446_;
  assign n3321_li = new_n3156_;
  assign n3324_li = new_n3158_;
  assign n3327_li = new_n3160_;
  assign n3330_li = new_n2448_;
  assign n3333_li = new_n3164_;
  assign n3336_li = new_n3166_;
  assign n3339_li = new_n3168_;
  assign n3342_li = new_n2450_;
  assign n3345_li = new_n3172_;
  assign n3348_li = new_n3174_;
  assign n3351_li = new_n3176_;
  assign n3354_li = new_n2452_;
  assign n3357_li = new_n3180_;
  assign n3360_li = new_n3182_;
  assign n3363_li = new_n3184_;
  assign n3366_li = new_n2454_;
  assign n3369_li = new_n3188_;
  assign n3372_li = new_n3190_;
  assign n3375_li = new_n3192_;
  assign n3378_li = new_n2456_;
  assign n3381_li = new_n3196_;
  assign n3384_li = new_n3198_;
  assign n3387_li = new_n3200_;
  assign n3390_li = new_n2458_;
  assign n3393_li = new_n3204_;
  assign n3396_li = new_n3206_;
  assign n3399_li = new_n3208_;
  assign n3402_li = new_n2460_;
  assign n3405_li = new_n3212_;
  assign n3408_li = new_n3214_;
  assign n3411_li = new_n3216_;
  assign n3414_li = new_n2462_;
  assign n3417_li = new_n3220_;
  assign n3420_li = new_n3222_;
  assign n3423_li = new_n3224_;
  assign n3426_li = new_n2464_;
  assign n3429_li = new_n3228_;
  assign n3432_li = new_n3230_;
  assign n3435_li = new_n3232_;
  assign n3438_li = new_n2466_;
  assign n3441_li = new_n3236_;
  assign n3444_li = new_n3238_;
  assign n3447_li = new_n3240_;
  assign n3450_li = new_n2468_;
  assign n3453_li = new_n3244_;
  assign n3456_li = new_n3246_;
  assign n3459_li = new_n3248_;
  assign n3462_li = new_n2470_;
  assign n3465_li = new_n3252_;
  assign n3468_li = new_n3254_;
  assign n3471_li = new_n3256_;
  assign n3474_li = new_n2472_;
  assign n3477_li = new_n3260_;
  assign n3480_li = new_n3262_;
  assign n3483_li = new_n3264_;
  assign n3486_li = new_n2474_;
  assign n3489_li = new_n3268_;
  assign n3492_li = new_n3270_;
  assign n3495_li = new_n3272_;
  assign n3498_li = new_n2476_;
  assign n3501_li = new_n3276_;
  assign n3504_li = new_n3278_;
  assign n3507_li = new_n3280_;
  assign n3510_li = new_n2478_;
  assign n3513_li = new_n3284_;
  assign n3516_li = new_n3286_;
  assign n3519_li = new_n3288_;
  assign n3522_li = new_n2480_;
  assign n3525_li = new_n3292_;
  assign n3528_li = new_n3294_;
  assign n3531_li = new_n3296_;
  assign n3534_li = new_n2482_;
  assign n3537_li = new_n3300_;
  assign n3540_li = new_n3302_;
  assign n3543_li = new_n3304_;
  assign n3546_li = new_n2484_;
  assign n3549_li = new_n3308_;
  assign n3552_li = new_n3310_;
  assign n3555_li = new_n3312_;
  assign n3558_li = new_n2486_;
  assign n3561_li = new_n3316_;
  assign n3564_li = new_n3318_;
  assign n3567_li = new_n3320_;
  assign n3570_li = new_n2488_;
  assign n3573_li = new_n3324_;
  assign n3576_li = new_n3326_;
  assign n3579_li = new_n3328_;
  assign n3582_li = new_n2490_;
  assign n3585_li = new_n3332_;
  assign n3588_li = new_n3334_;
  assign n3591_li = new_n3336_;
  assign n3594_li = new_n2492_;
  assign n3597_li = new_n3340_;
  assign n3600_li = new_n3342_;
  assign n3603_li = new_n3344_;
  assign n3606_li = new_n2494_;
  assign n3609_li = new_n3348_;
  assign n3612_li = new_n3350_;
  assign n3615_li = new_n3352_;
  assign n3618_li = new_n2496_;
  assign n3621_li = new_n3356_;
  assign n3624_li = new_n3358_;
  assign n3627_li = new_n3360_;
  assign n3630_li = new_n2498_;
  assign n3633_li = new_n3364_;
  assign n3636_li = new_n3366_;
  assign n3639_li = new_n3368_;
  assign n3642_li = new_n2500_;
  assign n3645_li = new_n3372_;
  assign n3648_li = new_n3374_;
  assign n3651_li = new_n3376_;
  assign n3654_li = new_n2502_;
  assign n3657_li = new_n3380_;
  assign n3666_li = new_n2504_;
  assign n3669_li = new_n3384_;
  assign n3678_li = new_n2506_;
  assign n3687_li = new_n10128_;
  assign n3690_li = new_n2508_;
  assign n3702_li = new_n2510_;
  assign n3711_li = new_n10117_;
  assign n3714_li = new_n2512_;
  assign n3726_li = new_n2514_;
  assign n3735_li = new_n10095_;
  assign n3738_li = new_n2516_;
  assign n3750_li = new_n2518_;
  assign n3753_li = new_n3406_;
  assign n3759_li = new_n10033_;
  assign n3762_li = new_n2520_;
  assign n3765_li = new_n3412_;
  assign n3774_li = new_n2522_;
  assign n3777_li = new_n3416_;
  assign n3786_li = new_n2524_;
  assign n3789_li = new_n3420_;
  assign n3792_li = new_n3422_;
  assign n3795_li = new_n3424_;
  assign n3798_li = new_n2526_;
  assign n3801_li = new_n3428_;
  assign n3810_li = new_n2528_;
  assign n3813_li = new_n3432_;
  assign n3822_li = new_n2530_;
  assign n3825_li = new_n3436_;
  assign n3834_li = new_n2532_;
  assign n3843_li = new_n10034_;
  assign n3846_li = new_n2534_;
  assign n3867_li = new_n9977_;
  assign n3891_li = new_n9976_;
  assign n3915_li = new_n9987_;
  assign n3930_li = new_n2548_;
  assign n3933_li = new_n3452_;
  assign n3936_li = new_n3454_;
  assign n3942_li = new_n2550_;
  assign n3945_li = new_n3458_;
  assign n3948_li = new_n3460_;
  assign n3954_li = new_n2552_;
  assign n3957_li = new_n3464_;
  assign n3963_li = new_n10161_;
  assign n3966_li = new_n2554_;
  assign n3969_li = new_n3470_;
  assign n3975_li = new_n4244_;
  assign n3978_li = new_n2556_;
  assign n3987_li = new_n10156_;
  assign n3990_li = new_n2558_;
  assign n4002_li = new_n2560_;
  assign n4011_li = new_n10147_;
  assign n4014_li = new_n2562_;
  assign n4026_li = new_n2564_;
  assign n4035_li = new_n10140_;
  assign n4038_li = new_n2566_;
  assign n4050_li = new_n2568_;
  assign n4053_li = new_n3494_;
  assign n4059_li = new_n10518_;
  assign n4062_li = new_n2570_;
  assign n4065_li = new_n3500_;
  assign n4098_li = new_n2576_;
  assign n4107_li = new_n3932_;
  assign n4119_li = new_n9990_;
  assign n4131_li = new_n3874_;
  assign n4143_li = new_n9989_;
  assign n4155_li = new_n3878_;
  assign n4167_li = new_n9696_;
  assign n4179_li = new_n3914_;
  assign n4182_li = new_n2590_;
  assign n4185_li = new_n3520_;
  assign n4188_li = new_n3522_;
  assign n4194_li = new_n2592_;
  assign n4197_li = new_n3526_;
  assign n4200_li = new_n3528_;
  assign n4206_li = new_n2594_;
  assign n4209_li = new_n3532_;
  assign n4212_li = new_n3534_;
  assign n4215_li = new_n3536_;
  assign n4227_li = new_n9933_;
  assign n4230_li = new_n2598_;
  assign n4233_li = new_n3542_;
  assign n4236_li = new_n3544_;
  assign n4239_li = new_n3546_;
  assign n4242_li = new_n2600_;
  assign n4251_li = new_n9939_;
  assign n4263_li = new_n9947_;
  assign n4275_li = new_n9955_;
  assign n4278_li = new_n2606_;
  assign n4287_li = new_n9728_;
  assign n4290_li = new_n2608_;
  assign n4293_li = new_n3562_;
  assign n4299_li = new_n9677_;
  assign n4302_li = new_n2610_;
  assign n4305_li = new_n3568_;
  assign n4311_li = new_n9553_;
  assign n4314_li = new_n2612_;
  assign n4323_li = new_n9763_;
  assign n4326_li = new_n2614_;
  assign n4335_li = new_n9736_;
  assign n4338_li = new_n2616_;
  assign n4347_li = new_n9775_;
  assign n4350_li = new_n2618_;
  assign n4359_li = new_n9911_;
  assign n4362_li = new_n2620_;
  assign n4365_li = new_n3590_;
  assign n4371_li = new_n9687_;
  assign n4374_li = new_n2622_;
  assign n4383_li = new_n9961_;
  assign n4395_li = new_n9968_;
  assign n4407_li = new_n9975_;
  assign n4410_li = new_n2628_;
  assign n4413_li = new_n3604_;
  assign n4416_li = new_n3606_;
  assign n4419_li = new_n3608_;
  assign n4422_li = new_n2630_;
  assign n4425_li = new_n3612_;
  assign n4428_li = new_n3614_;
  assign n4431_li = new_n3616_;
  assign n4434_li = new_n2632_;
  assign n4437_li = new_n3620_;
  assign n4440_li = new_n3622_;
  assign n4443_li = new_n3624_;
  assign n4446_li = new_n2634_;
  assign n4449_li = new_n3628_;
  assign n4452_li = new_n3630_;
  assign n4455_li = new_n3632_;
  assign n4458_li = new_n2636_;
  assign n4461_li = new_n3636_;
  assign n4464_li = new_n3638_;
  assign n4467_li = new_n3640_;
  assign n4470_li = new_n2638_;
  assign n4473_li = new_n3644_;
  assign n4476_li = new_n3646_;
  assign n4479_li = new_n3648_;
  assign n4482_li = new_n2640_;
  assign n4485_li = new_n3652_;
  assign n4488_li = new_n3654_;
  assign n4494_li = new_n2642_;
  assign n4497_li = new_n3658_;
  assign n4500_li = new_n3660_;
  assign n4503_li = new_n3662_;
  assign n4506_li = new_n2644_;
  assign n4509_li = new_n3666_;
  assign n4512_li = new_n3668_;
  assign n4515_li = new_n3670_;
  assign n4518_li = new_n2646_;
  assign n4521_li = new_n3674_;
  assign n4524_li = new_n3676_;
  assign n4527_li = new_n3678_;
  assign n4530_li = new_n2648_;
  assign n4533_li = new_n3682_;
  assign n4536_li = new_n3684_;
  assign n4539_li = new_n3686_;
  assign n4542_li = new_n2650_;
  assign n4545_li = new_n3690_;
  assign n4548_li = new_n3692_;
  assign n4554_li = new_n2652_;
  assign n4557_li = new_n3696_;
  assign n4560_li = new_n3698_;
  assign n4563_li = new_n3700_;
  assign n4566_li = new_n2654_;
  assign n4569_li = new_n3704_;
  assign n4572_li = new_n3706_;
  assign n4575_li = new_n3708_;
  assign n4578_li = new_n2656_;
  assign n4581_li = new_n3712_;
  assign n4584_li = new_n3714_;
  assign n4587_li = new_n3716_;
  assign n4590_li = new_n2658_;
  assign n4593_li = new_n3720_;
  assign n4596_li = new_n3722_;
  assign n4599_li = new_n3724_;
  assign n4602_li = new_n2660_;
  assign n4605_li = new_n3728_;
  assign n4608_li = new_n3730_;
  assign n4611_li = new_n3732_;
  assign n4614_li = new_n2662_;
  assign n4617_li = new_n3736_;
  assign n4620_li = new_n3738_;
  assign n4623_li = new_n3740_;
  assign n4626_li = new_n2664_;
  assign n4629_li = new_n3744_;
  assign n4632_li = new_n3746_;
  assign n4635_li = new_n3748_;
  assign n4638_li = new_n2666_;
  assign n4641_li = new_n3752_;
  assign n4644_li = new_n3754_;
  assign n4647_li = new_n3756_;
  assign n4650_li = new_n2668_;
  assign n4653_li = new_n3760_;
  assign n4656_li = new_n3762_;
  assign n4659_li = new_n3764_;
  assign n4662_li = new_n2670_;
  assign n4665_li = new_n3768_;
  assign n4668_li = new_n3770_;
  assign n4671_li = new_n3772_;
  assign n4674_li = new_n2672_;
  assign n4677_li = new_n3776_;
  assign n4680_li = new_n3778_;
  assign n4683_li = new_n3780_;
  assign n4686_li = new_n2674_;
  assign n4689_li = new_n3784_;
  assign n4692_li = new_n3786_;
  assign n4695_li = new_n3788_;
  assign n4698_li = new_n2676_;
  assign n4701_li = new_n3792_;
  assign n4704_li = new_n3794_;
  assign n4707_li = new_n3796_;
  assign n4710_li = new_n2678_;
  assign n4713_li = new_n3800_;
  assign n4716_li = new_n3802_;
  assign n4719_li = new_n3804_;
  assign n4722_li = new_n2680_;
  assign n4725_li = new_n3808_;
  assign n4728_li = new_n3810_;
  assign n4731_li = new_n3812_;
  assign n4734_li = new_n2682_;
  assign n4737_li = new_n3816_;
  assign n4740_li = new_n3818_;
  assign n4743_li = new_n3820_;
  assign n6382_i2 = new_n3996_;
  assign n6383_i2 = new_n3998_;
  assign n6419_i2 = new_n4008_;
  assign n6420_i2 = new_n4010_;
  assign n6435_i2 = new_n4018_;
  assign n6436_i2 = new_n4020_;
  assign n6448_i2 = new_n4024_;
  assign n6449_i2 = new_n4026_;
  assign n6613_i2 = new_n9845_;
  assign n6614_i2 = new_n9878_;
  assign n6641_i2 = new_n4060_;
  assign n6658_i2 = new_n4062_;
  assign n6757_i2 = new_n9674_;
  assign n6756_i2 = new_n9684_;
  assign n7116_i2 = new_n9901_;
  assign n7156_i2 = new_n10520_;
  assign n6549_i2 = new_n4032_;
  assign n6550_i2 = new_n4034_;
  assign n7357_i2 = new_n10063_;
  assign n7358_i2 = new_n9561_;
  assign n7359_i2 = new_n10076_;
  assign n7360_i2 = new_n9577_;
  assign n6621_i2 = new_n10522_;
  assign n6623_i2 = new_n10525_;
  assign n6625_i2 = new_n10528_;
  assign n6626_i2 = new_n4050_;
  assign n6627_i2 = new_n10531_;
  assign n6628_i2 = new_n4054_;
  assign n6629_i2 = new_n4056_;
  assign n6630_i2 = new_n4058_;
  assign n6669_i2 = new_n4064_;
  assign n7449_i2 = new_n10093_;
  assign n7450_i2 = new_n9593_;
  assign n7451_i2 = new_n9607_;
  assign n7452_i2 = new_n10112_;
  assign n6682_i2 = new_n4066_;
  assign n6683_i2 = new_n4068_;
  assign n6684_i2 = new_n4070_;
  assign n6685_i2 = new_n4072_;
  assign n7463_i2 = new_n9870_;
  assign n6686_i2 = new_n4074_;
  assign n6687_i2 = new_n4076_;
  assign n6688_i2 = new_n4078_;
  assign n6689_i2 = new_n4080_;
  assign n6772_i2 = new_n4090_;
  assign n6773_i2 = new_n4092_;
  assign n6774_i2 = new_n4094_;
  assign n6775_i2 = new_n4096_;
  assign G3467_i2 = new_n9844_;
  assign G2810_i2 = n7463_i2;
  assign n6833_i2 = new_n4102_;
  assign n6945_i2 = new_n10533_;
  assign n6947_i2 = new_n10366_;
  assign n6949_i2 = new_n10534_;
  assign n6951_i2 = new_n4132_;
  assign n6888_i2 = new_n4114_;
  assign n6889_i2 = new_n4116_;
  assign n6936_i2 = new_n4124_;
  assign n6954_i2 = new_n4138_;
  assign n6955_i2 = new_n10227_;
  assign n6956_i2 = new_n4142_;
  assign n6957_i2 = new_n10244_;
  assign n6958_i2 = new_n4146_;
  assign n6982_i2 = new_n10535_;
  assign n6984_i2 = new_n10536_;
  assign n6974_i2 = new_n4148_;
  assign n6975_i2 = new_n4150_;
  assign n6999_i2 = new_n10226_;
  assign n7015_i2 = new_n10359_;
  assign n7016_i2 = new_n4162_;
  assign n7017_i2 = new_n4164_;
  assign n7018_i2 = new_n4166_;
  assign n7005_i2 = new_n4158_;
  assign n7019_i2 = new_n4168_;
  assign n7022_i2 = new_n4170_;
  assign n7023_i2 = new_n4172_;
  assign n7132_i2 = new_n10280_;
  assign n7133_i2 = new_n10327_;
  assign n7135_i2 = new_n10326_;
  assign n7136_i2 = new_n10279_;
  assign n7175_i2 = new_n10537_;
  assign n7155_i2 = new_n10239_;
  assign G3060_i2 = new_n10134_;
  assign n7383_i2 = new_n9698_;
  assign G3802_i2 = new_n9857_;
  assign G3859_i2 = new_n9890_;
  assign n7355_i2 = new_n10261_;
  assign n7356_i2 = new_n10309_;
  assign G4054_i2 = new_n9849_;
  assign G4068_i2 = new_n9888_;
  assign n7384_i2 = new_n9697_;
  assign n7387_i2 = new_n4486_;
  assign n7388_i2 = new_n10256_;
  assign n7389_i2 = new_n10304_;
  assign n7386_i2 = new_n4484_;
  assign n7453_i2 = new_n4568_;
  assign n7431_i2 = new_n10213_;
  assign n7432_i2 = new_n10250_;
  assign n7433_i2 = new_n10294_;
  assign n7430_i2 = new_n10230_;
  assign n7485_i2 = new_n10267_;
  assign n7486_i2 = new_n10315_;
  assign G2508_i2 = new_n10201_;
  assign G2486_i2 = new_n10300_;
  assign n7245_i2 = new_n9719_;
  assign n7246_i2 = new_n9813_;
  assign n3756_lo_buf_i2 = new_n9708_;
  assign n4056_lo_buf_i2 = new_n9701_;
  assign G3474_i2 = new_n10249_;
  assign G2817_i2 = G2486_i2;
  assign n7396_i2 = new_n4492_;
  assign n7398_i2 = new_n4494_;
  assign n7400_i2 = new_n4496_;
  assign n7401_i2 = new_n4498_;
  assign n7402_i2 = new_n4500_;
  assign n7403_i2 = new_n4502_;
  assign n7404_i2 = new_n9714_;
  assign n7405_i2 = new_n9811_;
  assign G2711_i2 = new_n10270_;
  assign G2828_i2 = new_n10299_;
  assign n7490_i2 = new_n4620_;
  assign n7527_i2 = new_n9806_;
  assign n7528_i2 = new_n9749_;
  assign n7529_i2 = new_n9808_;
  assign n7530_i2 = new_n9751_;
  assign n7523_i2 = new_n9809_;
  assign n7524_i2 = new_n9752_;
  assign n7525_i2 = new_n9807_;
  assign n7526_i2 = new_n9750_;
  assign n4296_lo_buf_i2 = new_n9918_;
  assign n4368_lo_buf_i2 = new_n9922_;
  assign G2466_i2 = new_n9923_;
  assign G2404_i2 = new_n9919_;
  assign n7534_i2 = new_n9713_;
  assign n7535_i2 = new_n9717_;
  assign n7536_i2 = new_n9779_;
  assign n7533_i2 = new_n9783_;
  assign G1060_i2 = new_n9819_;
  assign G963_i2 = new_n9830_;
  assign G2448_i2 = new_n10451_;
  assign G2685_i2 = new_n9995_;
  assign G2679_i2 = new_n10002_;
  assign G2774_i2 = ~new_n10004_;
  assign G2780_i2 = ~new_n10013_;
  assign G2759_i2 = new_n10009_;
  assign G2737_i2 = new_n10398_;
  assign G2850_i2 = new_n10410_;
  assign G3393_i2 = new_n10001_;
  assign G3404_i2 = new_n9994_;
  assign G3559_i2 = new_n10024_;
  assign G2744_i2 = new_n10429_;
  assign n3708_lo_buf_i2 = new_n9831_;
  assign n3840_lo_buf_i2 = new_n9812_;
  assign n4008_lo_buf_i2 = new_n9820_;
  assign n4104_lo_buf_i2 = new_n9810_;
  assign G1821_i2 = new_n9818_;
  assign G1734_i2 = new_n9829_;
  assign G3517_i2 = new_n10397_;
  assign G3533_i2 = new_n10423_;
  assign G3629_i2 = new_n10408_;
  assign G3645_i2 = new_n10438_;
  assign G2857_i2 = new_n10452_;
  assign G2731_i2 = new_n10455_;
  assign G2844_i2 = new_n10458_;
  assign n3732_lo_buf_i2 = new_n9925_;
  assign n4032_lo_buf_i2 = new_n9924_;
  assign G3552_i2 = new_n10435_;
  assign G2271_i2 = new_n10343_;
  assign n4248_lo_buf_i2 = new_n10347_;
  assign n4332_lo_buf_i2 = new_n10351_;
  assign n4344_lo_buf_i2 = new_n10355_;
  assign n4380_lo_buf_i2 = new_n10341_;
  assign G2398_i2 = new_n10349_;
  assign G2480_i2 = new_n10357_;
  assign G2418_i2 = new_n10353_;
  assign G1455_i2 = new_n10130_;
  assign G1449_i2 = new_n10119_;
  assign G1452_i2 = new_n10097_;
  assign G1425_i2 = new_n10163_;
  assign G1428_i2 = new_n10158_;
  assign G1419_i2 = new_n10149_;
  assign G1422_i2 = new_n10142_;
  assign n4308_lo_buf_i2 = new_n3570_;
  assign G2675_i2 = new_n10029_;
  assign G3035_i2 = new_n9942_;
  assign G3026_i2 = new_n9950_;
  assign G3029_i2 = new_n9928_;
  assign G3032_i2 = new_n9936_;
  assign G2999_i2 = new_n9770_;
  assign G3002_i2 = new_n9906_;
  assign G2770_i2 = new_n10011_;
  assign G3008_i2 = G2770_i2;
  assign G2073_i2 = n7156_i2;
  assign G2752_i2 = new_n9872_;
  assign G3005_i2 = G2752_i2;
  assign G5108_i2 = new_n10538_;
  assign G5135_i2 = new_n10539_;
  assign G5111_i2 = new_n10540_;
  assign G5138_i2 = new_n10541_;
  assign G3415_i2 = new_n10026_;
  assign G3386_i2 = new_n10542_;
  assign G3570_i2 = new_n10022_;
  assign G2430_i2 = new_n10368_;
  assign G3495_i2 = new_n10379_;
  assign G3621_i2 = new_n10390_;
  assign n4284_lo_buf_i2 = new_n10207_;
  assign n4356_lo_buf_i2 = new_n10211_;
  assign G2472_i2 = new_n10209_;
  assign G2410_i2 = new_n10205_;
  assign n3960_lo_buf_i2 = new_n10393_;
  assign n3972_lo_buf_i2 = new_n10394_;
  assign G2865_i2 = G2857_i2;
  assign G970_i2 = new_n9914_;
  assign n3684_lo_buf_i2 = new_n10338_;
  assign n4080_lo_buf_i2 = new_n10493_;
  assign n4092_lo_buf_i2 = new_n10503_;
  assign G1053_i2 = new_n10495_;
  assign G956_i2 = new_n10504_;
  assign G1147_i2 = n4059_li;
  assign G2705_i2 = new_n6554_;
  assign G2693_i2 = new_n6555_;
  assign G2696_i2 = new_n6556_;
  assign G2700_i2 = new_n6557_;
  assign G2915_i2 = new_n6558_;
  assign G2966_i2 = new_n6559_;
  assign G2540_i2 = new_n6560_;
  assign G2788_i2 = new_n6561_;
  assign G2792_i2 = new_n6562_;
  assign G2797_i2 = new_n10021_;
  assign G2804_i2 = G2797_i2;
  assign G1038_i2 = n6621_i2;
  assign G1044_i2 = n6623_i2;
  assign G1090_i2 = n6625_i2;
  assign G1096_i2 = n6627_i2;
  assign G1029_i2 = new_n10367_;
  assign G3942_i2 = n7388_i2;
  assign G3954_i2 = new_n10258_;
  assign G4011_i2 = n7389_i2;
  assign G4017_i2 = new_n10306_;
  assign G1141_i2 = new_n9710_;
  assign G1081_i2 = new_n9703_;
  assign G2146_i2 = new_n6563_;
  assign G2145_i2 = new_n6564_;
  assign G2144_i2 = new_n6565_;
  assign G2143_i2 = new_n6566_;
  assign G2142_i2 = new_n6567_;
  assign G2141_i2 = new_n6568_;
  assign G2140_i2 = new_n6569_;
  assign G2139_i2 = new_n6570_;
  assign G3769_i2 = new_n10030_;
  assign G3773_i2 = new_n9996_;
  assign G3768_i2 = new_n10028_;
  assign G4101_i2 = new_n6574_;
  assign G3161_i2 = ~new_n10031_;
  assign G4143_i2 = ~new_n6577_;
  assign G3828_i2 = ~new_n10032_;
  assign G3831_i2 = ~new_n10014_;
  assign G3334_i2 = new_n6579_;
  assign G3335_i2 = new_n6580_;
  assign G3180_i2 = new_n6584_;
  assign G3340_i2 = new_n6585_;
  assign G3339_i2 = new_n6586_;
  assign G3341_i2 = new_n6587_;
  assign G3234_i2 = new_n10012_;
  assign G3829_i2 = new_n6589_;
  assign G3338_i2 = new_n6590_;
  assign G3336_i2 = new_n6591_;
  assign G3770_i2 = new_n6593_;
  assign G3918_i2 = G3393_i2;
  assign G3774_i2 = new_n10027_;
  assign G3921_i2 = G3404_i2;
  assign G3832_i2 = new_n10025_;
  assign G3993_i2 = new_n10023_;
  assign G2076_i2 = G1455_i2;
  assign G2071_i2 = G1449_i2;
  assign G2072_i2 = G1452_i2;
  assign G2069_i2 = G1425_i2;
  assign G2070_i2 = G1428_i2;
  assign G2067_i2 = G1419_i2;
  assign G2068_i2 = G1422_i2;
  assign G4095_i2 = new_n6595_;
  assign G3272_i2 = G3035_i2;
  assign G3269_i2 = G3026_i2;
  assign G3270_i2 = G3029_i2;
  assign G3271_i2 = G3032_i2;
  assign G3265_i2 = G2999_i2;
  assign G3266_i2 = G3002_i2;
  assign G4137_i2 = new_n6597_;
  assign G3268_i2 = G3234_i2;
  assign G2361_i2 = new_n10519_;
  assign G3228_i2 = new_n9873_;
  assign G3267_i2 = G3228_i2;
  assign G2336_i2 = new_n6600_;
  assign G3459_i2 = new_n6603_;
  assign G3428_i2 = new_n6606_;
  assign G3438_i2 = new_n6609_;
  assign G3449_i2 = new_n6612_;
  assign G3421_i2 = new_n6615_;
  assign G3576_i2 = new_n6618_;
  assign G3303_i2 = new_n6621_;
  assign G3583_i2 = new_n6624_;
  assign G3594_i2 = new_n6627_;
  assign G3674_i2 = new_n6630_;
  assign G3685_i2 = new_n6639_;
  assign G4504_i2 = new_n6714_;
  assign G4180_i2 = new_n6781_;
  assign G5123_i2 = G5108_i2;
  assign G5142_i2 = G5135_i2;
  assign G5126_i2 = G5111_i2;
  assign G5144_i2 = G5138_i2;
  assign G3912_i2 = G3386_i2;
  assign G4417_i2 = new_n6888_;
  assign G4420_i2 = new_n6969_;
  assign G3969_i2 = new_n10381_;
  assign G4023_i2 = new_n10392_;
  assign G2720_i2 = new_n10486_;
  assign G2837_i2 = new_n10488_;
  assign G836_i2 = new_n10543_;
  assign G848_i2 = G836_i2;
  assign G813_i2 = new_n10544_;
  assign G825_i2 = G813_i2;
  assign G1876_i2 = new_n9913_;
  assign G4996_i2 = new_n10545_;
  assign G4984_i2 = new_n10546_;
  assign G4920_i2 = new_n10547_;
  assign G4923_i2 = new_n10548_;
  assign G4930_i2 = new_n10549_;
  assign G4933_i2 = new_n10550_;
  assign n4320_lo_buf_i2 = new_n10552_;
  assign G2424_i2 = new_n10554_;
  assign G3317_i2 = new_n7130_;
  assign G3503_i2 = new_n10407_;
  assign G3485_i2 = new_n10473_;
  assign G3611_i2 = new_n10476_;
  assign n3864_lo_buf_i2 = new_n10505_;
  assign n3888_lo_buf_i2 = new_n10508_;
  assign n4116_lo_buf_i2 = new_n10491_;
  assign n4128_lo_buf_i2 = new_n10496_;
  assign n4140_lo_buf_i2 = new_n10498_;
  assign n4152_lo_buf_i2 = new_n10499_;
  assign G1815_i2 = G1053_i2;
  assign G1728_i2 = G956_i2;
  assign G1035_i2 = new_n10523_;
  assign G1041_i2 = new_n10526_;
  assign G1087_i2 = new_n10529_;
  assign G1093_i2 = new_n10532_;
  assign G1132_i2 = n6945_i2;
  assign G1108_i2 = n6949_i2;
  assign G1138_i2 = n6982_i2;
  assign G1114_i2 = n6984_i2;
  assign G1807_i2 = new_n7141_;
  assign G2108_i2 = new_n7143_;
  assign G1126_i2 = n7175_i2;
  assign G1899_i2 = new_n7145_;
  assign G2134_i2 = new_n7147_;
  assign G1852_i2 = new_n7149_;
  assign G2116_i2 = new_n7151_;
  assign G2543_i2 = ~new_n10483_;
  assign G2727_i2 = new_n10479_;
  assign G2715_i2 = new_n10487_;
  assign G2832_i2 = new_n10489_;
  assign G1873_i2 = new_n9915_;
  assign G3291_i2 = new_n7156_;
  assign G5025_i2 = new_n7172_;
  assign G5036_i2 = new_n7188_;
  assign G3132_i2 = ~new_n7189_;
  assign G5038_i2 = new_n7190_;
  assign G5039_i2 = new_n7191_;
  assign G1150_i2 = new_n10555_;
  assign G1162_i2 = G1150_i2;
  assign G804_i2 = new_n10556_;
  assign G1172_i2 = G804_i2;
  assign n3984_lo_buf_i2 = new_n10434_;
  assign G1802_i2 = G1035_i2;
  assign G1804_i2 = G1041_i2;
  assign G1849_i2 = G1087_i2;
  assign G1851_i2 = G1093_i2;
  assign G2492_i2 = new_n7194_;
  assign G1799_i2 = G1029_i2;
  assign G4231_i2 = G3954_i2;
  assign G4234_i2 = new_n10257_;
  assign G4245_i2 = G4017_i2;
  assign G4247_i2 = new_n10305_;
  assign G1894_i2 = G1141_i2;
  assign G1846_i2 = G1081_i2;
  assign G4238_i2 = G3969_i2;
  assign G4249_i2 = G4023_i2;
  assign G2293_i2 = G1873_i2;
  assign G5022_i2 = G4996_i2;
  assign G5006_i2 = G4984_i2;
  assign G4944_i2 = G4920_i2;
  assign G4946_i2 = G4923_i2;
  assign G4954_i2 = G4930_i2;
  assign G4956_i2 = G4933_i2;
  assign G3546_i2 = new_n10472_;
  assign G3658_i2 = new_n10475_;
  assign G1344_i2 = n4320_lo_buf_i2;
  assign G2921_i2 = G2424_i2;
  assign n3912_lo_buf_i2 = new_n10509_;
  assign G1835_i2 = new_n7201_;
  assign G3810_i2 = new_n10480_;
  assign G3866_i2 = ~new_n10484_;
  assign G3811_i2 = new_n10481_;
  assign G2269_i2 = new_n7213_;
  assign G3812_i2 = new_n7217_;
  assign G3867_i2 = ~new_n10485_;
  assign G3868_i2 = ~new_n7225_;
  assign G3809_i2 = new_n10478_;
  assign G3716_i2 = ~new_n10482_;
  assign G4529_i2 = ~new_n7239_;
  assign G4670_i2 = new_n7259_;
  assign G4493_i2 = new_n7260_;
  assign G4580_i2 = new_n7261_;
  assign G3822_i2 = new_n7262_;
  assign G3877_i2 = new_n7263_;
  assign G4131_i2 = new_n7266_;
  assign G4170_i2 = ~new_n7269_;
  assign G4051_i2 = new_n7271_;
  assign G4065_i2 = new_n7273_;
  assign G4697_i2 = new_n7282_;
  assign G4706_i2 = new_n7291_;
  assign G2460_i2 = new_n10557_;
  assign G2454_i2 = new_n10558_;
  assign G2392_i2 = new_n10559_;
  assign G2386_i2 = new_n10560_;
  assign n4260_lo_buf_i2 = new_n10561_;
  assign n4272_lo_buf_i2 = new_n10562_;
  assign n4392_lo_buf_i2 = new_n10563_;
  assign n4404_lo_buf_i2 = new_n10564_;
  assign G1512_i2 = new_n10551_;
  assign G3135_i2 = new_n10553_;
  assign G2379_i2 = new_n7306_;
  assign n4164_lo_buf_i2 = new_n2586_;
  assign n4176_lo_buf_i2 = new_n2588_;
  assign n4224_lo_buf_i2 = new_n2596_;
  assign G2975_i2 = G2460_i2;
  assign G2978_i2 = G2454_i2;
  assign G2933_i2 = G2392_i2;
  assign G2936_i2 = G2386_i2;
  assign G1356_i2 = n4260_lo_buf_i2;
  assign G1359_i2 = n4272_lo_buf_i2;
  assign G1398_i2 = n4392_lo_buf_i2;
  assign G1401_i2 = n4404_lo_buf_i2;
  assign new_n8443_ = new_n3210_;
  assign new_n8444_ = new_n2690_;
  assign new_n8445_ = new_n3719_;
  assign new_n8446_ = new_n2771_;
  assign new_n8447_ = new_n3635_;
  assign new_n8448_ = new_n3549_;
  assign new_n8449_ = new_n4717_;
  assign new_n8450_ = new_n8449_;
  assign new_n8451_ = new_n8450_;
  assign new_n8452_ = new_n8451_;
  assign new_n8453_ = new_n8451_;
  assign new_n8454_ = new_n8450_;
  assign new_n8455_ = new_n8454_;
  assign new_n8456_ = new_n8454_;
  assign new_n8457_ = new_n8449_;
  assign new_n8458_ = new_n8457_;
  assign new_n8459_ = new_n8458_;
  assign new_n8460_ = new_n8457_;
  assign new_n8461_ = new_n3703_;
  assign new_n8462_ = new_n8461_;
  assign new_n8463_ = new_n8462_;
  assign new_n8464_ = new_n8462_;
  assign new_n8465_ = new_n8461_;
  assign new_n8466_ = new_n8465_;
  assign new_n8467_ = new_n8465_;
  assign new_n8468_ = new_n3702_;
  assign new_n8469_ = new_n8468_;
  assign new_n8470_ = new_n8469_;
  assign new_n8471_ = new_n8469_;
  assign new_n8472_ = new_n8468_;
  assign new_n8473_ = new_n8472_;
  assign new_n8474_ = new_n8472_;
  assign new_n8475_ = new_n2939_;
  assign new_n8476_ = new_n4716_;
  assign new_n8477_ = new_n4735_;
  assign new_n8478_ = new_n8477_;
  assign new_n8479_ = new_n8477_;
  assign new_n8480_ = new_n4736_;
  assign new_n8481_ = new_n8480_;
  assign new_n8482_ = new_n8480_;
  assign new_n8483_ = new_n3211_;
  assign new_n8484_ = new_n8483_;
  assign new_n8485_ = new_n8484_;
  assign new_n8486_ = new_n8483_;
  assign new_n8487_ = new_n3860_;
  assign new_n8488_ = new_n8487_;
  assign new_n8489_ = new_n3589_;
  assign new_n8490_ = new_n3490_;
  assign new_n8491_ = new_n3864_;
  assign new_n8492_ = new_n8491_;
  assign new_n8493_ = new_n3491_;
  assign new_n8494_ = new_n3887_;
  assign new_n8495_ = new_n8494_;
  assign new_n8496_ = new_n3893_;
  assign new_n8497_ = new_n8496_;
  assign new_n8498_ = new_n3585_;
  assign new_n8499_ = new_n3484_;
  assign new_n8500_ = new_n3485_;
  assign new_n8501_ = new_n3469_;
  assign new_n8502_ = new_n8501_;
  assign new_n8503_ = new_n3468_;
  assign new_n8504_ = new_n4784_;
  assign new_n8505_ = new_n4774_;
  assign new_n8506_ = new_n4787_;
  assign new_n8507_ = new_n3750_;
  assign new_n8508_ = new_n8507_;
  assign new_n8509_ = new_n8508_;
  assign new_n8510_ = new_n8509_;
  assign new_n8511_ = new_n8509_;
  assign new_n8512_ = new_n8508_;
  assign new_n8513_ = new_n8512_;
  assign new_n8514_ = new_n8512_;
  assign new_n8515_ = new_n8507_;
  assign new_n8516_ = new_n8515_;
  assign new_n8517_ = new_n8515_;
  assign new_n8518_ = new_n3603_;
  assign new_n8519_ = new_n3512_;
  assign new_n8520_ = new_n3742_;
  assign new_n8521_ = new_n8520_;
  assign new_n8522_ = new_n8521_;
  assign new_n8523_ = new_n8522_;
  assign new_n8524_ = new_n8522_;
  assign new_n8525_ = new_n8521_;
  assign new_n8526_ = new_n8525_;
  assign new_n8527_ = new_n8520_;
  assign new_n8528_ = new_n8527_;
  assign new_n8529_ = new_n8527_;
  assign new_n8530_ = new_n3513_;
  assign new_n8531_ = new_n3727_;
  assign new_n8532_ = new_n8531_;
  assign new_n8533_ = new_n8532_;
  assign new_n8534_ = new_n8533_;
  assign new_n8535_ = new_n8533_;
  assign new_n8536_ = new_n8532_;
  assign new_n8537_ = new_n8536_;
  assign new_n8538_ = new_n8536_;
  assign new_n8539_ = new_n8531_;
  assign new_n8540_ = new_n8539_;
  assign new_n8541_ = new_n8539_;
  assign new_n8542_ = new_n3735_;
  assign new_n8543_ = new_n8542_;
  assign new_n8544_ = new_n8543_;
  assign new_n8545_ = new_n8544_;
  assign new_n8546_ = new_n8544_;
  assign new_n8547_ = new_n8543_;
  assign new_n8548_ = new_n8547_;
  assign new_n8549_ = new_n8542_;
  assign new_n8550_ = new_n8549_;
  assign new_n8551_ = new_n8549_;
  assign new_n8552_ = new_n3601_;
  assign new_n8553_ = new_n3508_;
  assign new_n8554_ = new_n3509_;
  assign new_n8555_ = new_n3595_;
  assign new_n8556_ = new_n8555_;
  assign new_n8557_ = new_n3498_;
  assign new_n8558_ = new_n3499_;
  assign new_n8559_ = new_n3594_;
  assign new_n8560_ = new_n4816_;
  assign new_n8561_ = new_n4806_;
  assign new_n8562_ = new_n4819_;
  assign new_n8563_ = new_n4829_;
  assign new_n8564_ = new_n3567_;
  assign new_n8565_ = new_n8564_;
  assign new_n8566_ = new_n3410_;
  assign new_n8567_ = new_n3411_;
  assign new_n8568_ = new_n3566_;
  assign new_n8569_ = new_n3561_;
  assign new_n8570_ = new_n3402_;
  assign new_n8571_ = new_n3403_;
  assign new_n8572_ = new_n3581_;
  assign new_n8573_ = new_n3396_;
  assign new_n8574_ = new_n3397_;
  assign new_n8575_ = new_n3577_;
  assign new_n8576_ = new_n3390_;
  assign new_n8577_ = new_n3391_;
  assign new_n8578_ = new_n4854_;
  assign new_n8579_ = new_n4844_;
  assign new_n8580_ = new_n4864_;
  assign new_n8581_ = new_n4874_;
  assign new_n8582_ = new_n3541_;
  assign new_n8583_ = new_n3450_;
  assign new_n8584_ = new_n3451_;
  assign new_n8585_ = new_n3557_;
  assign new_n8586_ = new_n3448_;
  assign new_n8587_ = new_n3449_;
  assign new_n8588_ = new_n3555_;
  assign new_n8589_ = new_n3446_;
  assign new_n8590_ = new_n3447_;
  assign new_n8591_ = new_n3553_;
  assign new_n8592_ = new_n3442_;
  assign new_n8593_ = new_n3443_;
  assign new_n8594_ = new_n4897_;
  assign new_n8595_ = new_n4887_;
  assign new_n8596_ = new_n4907_;
  assign new_n8597_ = new_n4917_;
  assign new_n8598_ = new_n3829_;
  assign new_n8599_ = new_n3841_;
  assign new_n8600_ = new_n8599_;
  assign new_n8601_ = new_n3921_;
  assign new_n8602_ = new_n8601_;
  assign new_n8603_ = new_n8601_;
  assign new_n8604_ = new_n4925_;
  assign new_n8605_ = new_n4227_;
  assign new_n8606_ = new_n4112_;
  assign new_n8607_ = new_n8606_;
  assign new_n8608_ = new_n8606_;
  assign new_n8609_ = new_n4123_;
  assign new_n8610_ = new_n8609_;
  assign new_n8611_ = new_n4210_;
  assign new_n8612_ = new_n8611_;
  assign new_n8613_ = new_n8612_;
  assign new_n8614_ = new_n8612_;
  assign new_n8615_ = new_n8611_;
  assign new_n8616_ = new_n4422_;
  assign new_n8617_ = new_n8616_;
  assign new_n8618_ = new_n8617_;
  assign new_n8619_ = new_n8618_;
  assign new_n8620_ = new_n8617_;
  assign new_n8621_ = new_n8616_;
  assign new_n8622_ = new_n8621_;
  assign new_n8623_ = new_n8621_;
  assign new_n8624_ = new_n4281_;
  assign new_n8625_ = new_n8624_;
  assign new_n8626_ = new_n4423_;
  assign new_n8627_ = new_n8626_;
  assign new_n8628_ = new_n8627_;
  assign new_n8629_ = new_n8628_;
  assign new_n8630_ = new_n8627_;
  assign new_n8631_ = new_n8626_;
  assign new_n8632_ = new_n8631_;
  assign new_n8633_ = new_n8631_;
  assign new_n8634_ = new_n4280_;
  assign new_n8635_ = new_n8634_;
  assign new_n8636_ = new_n4424_;
  assign new_n8637_ = new_n8636_;
  assign new_n8638_ = new_n8637_;
  assign new_n8639_ = new_n8637_;
  assign new_n8640_ = new_n8636_;
  assign new_n8641_ = new_n4425_;
  assign new_n8642_ = new_n8641_;
  assign new_n8643_ = new_n8642_;
  assign new_n8644_ = new_n8642_;
  assign new_n8645_ = new_n8641_;
  assign new_n8646_ = new_n4420_;
  assign new_n8647_ = new_n8646_;
  assign new_n8648_ = new_n8647_;
  assign new_n8649_ = new_n8647_;
  assign new_n8650_ = new_n8646_;
  assign new_n8651_ = new_n4421_;
  assign new_n8652_ = new_n8651_;
  assign new_n8653_ = new_n8652_;
  assign new_n8654_ = new_n8652_;
  assign new_n8655_ = new_n8651_;
  assign new_n8656_ = new_n4426_;
  assign new_n8657_ = new_n8656_;
  assign new_n8658_ = new_n8657_;
  assign new_n8659_ = new_n8657_;
  assign new_n8660_ = new_n8656_;
  assign new_n8661_ = new_n4427_;
  assign new_n8662_ = new_n8661_;
  assign new_n8663_ = new_n8662_;
  assign new_n8664_ = new_n8662_;
  assign new_n8665_ = new_n8661_;
  assign new_n8666_ = new_n4937_;
  assign new_n8667_ = new_n4929_;
  assign new_n8668_ = new_n3831_;
  assign new_n8669_ = new_n3842_;
  assign new_n8670_ = new_n8669_;
  assign new_n8671_ = new_n3922_;
  assign new_n8672_ = new_n8671_;
  assign new_n8673_ = new_n8671_;
  assign new_n8674_ = new_n4941_;
  assign new_n8675_ = new_n4223_;
  assign new_n8676_ = new_n4119_;
  assign new_n8677_ = new_n8676_;
  assign new_n8678_ = new_n8676_;
  assign new_n8679_ = new_n4121_;
  assign new_n8680_ = new_n8679_;
  assign new_n8681_ = new_n4225_;
  assign new_n8682_ = new_n8681_;
  assign new_n8683_ = new_n8682_;
  assign new_n8684_ = new_n8681_;
  assign new_n8685_ = new_n4412_;
  assign new_n8686_ = new_n8685_;
  assign new_n8687_ = new_n8686_;
  assign new_n8688_ = new_n8687_;
  assign new_n8689_ = new_n8686_;
  assign new_n8690_ = new_n8685_;
  assign new_n8691_ = new_n8690_;
  assign new_n8692_ = new_n8690_;
  assign new_n8693_ = new_n4410_;
  assign new_n8694_ = new_n8693_;
  assign new_n8695_ = new_n4413_;
  assign new_n8696_ = new_n8695_;
  assign new_n8697_ = new_n8696_;
  assign new_n8698_ = new_n8697_;
  assign new_n8699_ = new_n8696_;
  assign new_n8700_ = new_n8695_;
  assign new_n8701_ = new_n8700_;
  assign new_n8702_ = new_n8700_;
  assign new_n8703_ = new_n4411_;
  assign new_n8704_ = new_n8703_;
  assign new_n8705_ = new_n4414_;
  assign new_n8706_ = new_n8705_;
  assign new_n8707_ = new_n8706_;
  assign new_n8708_ = new_n8706_;
  assign new_n8709_ = new_n8705_;
  assign new_n8710_ = new_n4415_;
  assign new_n8711_ = new_n8710_;
  assign new_n8712_ = new_n8711_;
  assign new_n8713_ = new_n8711_;
  assign new_n8714_ = new_n8710_;
  assign new_n8715_ = new_n4418_;
  assign new_n8716_ = new_n8715_;
  assign new_n8717_ = new_n8716_;
  assign new_n8718_ = new_n8716_;
  assign new_n8719_ = new_n8715_;
  assign new_n8720_ = new_n4419_;
  assign new_n8721_ = new_n8720_;
  assign new_n8722_ = new_n8721_;
  assign new_n8723_ = new_n8721_;
  assign new_n8724_ = new_n8720_;
  assign new_n8725_ = new_n4416_;
  assign new_n8726_ = new_n8725_;
  assign new_n8727_ = new_n8726_;
  assign new_n8728_ = new_n8726_;
  assign new_n8729_ = new_n8725_;
  assign new_n8730_ = new_n4417_;
  assign new_n8731_ = new_n8730_;
  assign new_n8732_ = new_n8731_;
  assign new_n8733_ = new_n8731_;
  assign new_n8734_ = new_n8730_;
  assign new_n8735_ = new_n4953_;
  assign new_n8736_ = new_n4945_;
  assign new_n8737_ = new_n4965_;
  assign new_n8738_ = new_n4960_;
  assign new_n8739_ = new_n4966_;
  assign new_n8740_ = new_n4959_;
  assign new_n8741_ = new_n4975_;
  assign new_n8742_ = new_n8741_;
  assign new_n8743_ = new_n8741_;
  assign new_n8744_ = new_n4974_;
  assign new_n8745_ = new_n8744_;
  assign new_n8746_ = new_n8744_;
  assign new_n8747_ = new_n4976_;
  assign new_n8748_ = new_n8747_;
  assign new_n8749_ = new_n8747_;
  assign new_n8750_ = new_n4973_;
  assign new_n8751_ = new_n8750_;
  assign new_n8752_ = new_n8750_;
  assign new_n8753_ = new_n4261_;
  assign new_n8754_ = new_n8753_;
  assign new_n8755_ = new_n8753_;
  assign new_n8756_ = new_n4260_;
  assign new_n8757_ = new_n8756_;
  assign new_n8758_ = new_n8756_;
  assign new_n8759_ = new_n5012_;
  assign new_n8760_ = new_n5007_;
  assign new_n8761_ = new_n5013_;
  assign new_n8762_ = new_n5006_;
  assign new_n8763_ = new_n5022_;
  assign new_n8764_ = new_n8763_;
  assign new_n8765_ = new_n8763_;
  assign new_n8766_ = new_n5021_;
  assign new_n8767_ = new_n8766_;
  assign new_n8768_ = new_n8766_;
  assign new_n8769_ = new_n5023_;
  assign new_n8770_ = new_n8769_;
  assign new_n8771_ = new_n8769_;
  assign new_n8772_ = new_n5020_;
  assign new_n8773_ = new_n8772_;
  assign new_n8774_ = new_n8772_;
  assign new_n8775_ = new_n4408_;
  assign new_n8776_ = new_n8775_;
  assign new_n8777_ = new_n8775_;
  assign new_n8778_ = new_n4409_;
  assign new_n8779_ = new_n8778_;
  assign new_n8780_ = new_n8778_;
  assign new_n8781_ = new_n3573_;
  assign new_n8782_ = new_n8781_;
  assign new_n8783_ = new_n5049_;
  assign new_n8784_ = new_n4204_;
  assign new_n8785_ = new_n4109_;
  assign new_n8786_ = new_n4111_;
  assign new_n8787_ = new_n3903_;
  assign new_n8788_ = new_n8787_;
  assign new_n8789_ = new_n8787_;
  assign new_n8790_ = new_n4274_;
  assign new_n8791_ = new_n4275_;
  assign new_n8792_ = new_n4276_;
  assign new_n8793_ = new_n8792_;
  assign new_n8794_ = new_n4277_;
  assign new_n8795_ = new_n8794_;
  assign new_n8796_ = new_n4278_;
  assign new_n8797_ = new_n8796_;
  assign new_n8798_ = new_n4279_;
  assign new_n8799_ = new_n8798_;
  assign new_n8800_ = new_n5084_;
  assign new_n8801_ = new_n5085_;
  assign new_n8802_ = new_n4283_;
  assign new_n8803_ = new_n8802_;
  assign new_n8804_ = new_n8802_;
  assign new_n8805_ = new_n4282_;
  assign new_n8806_ = new_n8805_;
  assign new_n8807_ = new_n8805_;
  assign new_n8808_ = new_n5098_;
  assign new_n8809_ = new_n4191_;
  assign new_n8810_ = new_n4107_;
  assign new_n8811_ = new_n4105_;
  assign new_n8812_ = new_n4264_;
  assign new_n8813_ = new_n4265_;
  assign new_n8814_ = new_n4266_;
  assign new_n8815_ = new_n8814_;
  assign new_n8816_ = new_n4267_;
  assign new_n8817_ = new_n8816_;
  assign new_n8818_ = new_n4268_;
  assign new_n8819_ = new_n8818_;
  assign new_n8820_ = new_n4269_;
  assign new_n8821_ = new_n8820_;
  assign new_n8822_ = new_n5125_;
  assign new_n8823_ = new_n5126_;
  assign new_n8824_ = new_n4262_;
  assign new_n8825_ = new_n8824_;
  assign new_n8826_ = new_n8824_;
  assign new_n8827_ = new_n4263_;
  assign new_n8828_ = new_n8827_;
  assign new_n8829_ = new_n8827_;
  assign new_n8830_ = new_n5139_;
  assign new_n8831_ = new_n3862_;
  assign new_n8832_ = new_n3866_;
  assign new_n8833_ = new_n3806_;
  assign new_n8834_ = new_n8833_;
  assign new_n8835_ = new_n8834_;
  assign new_n8836_ = new_n8835_;
  assign new_n8837_ = new_n8836_;
  assign new_n8838_ = new_n8837_;
  assign new_n8839_ = new_n8837_;
  assign new_n8840_ = new_n8836_;
  assign new_n8841_ = new_n8840_;
  assign new_n8842_ = new_n8840_;
  assign new_n8843_ = new_n8835_;
  assign new_n8844_ = new_n8843_;
  assign new_n8845_ = new_n8844_;
  assign new_n8846_ = new_n8844_;
  assign new_n8847_ = new_n8843_;
  assign new_n8848_ = new_n8847_;
  assign new_n8849_ = new_n8847_;
  assign new_n8850_ = new_n8834_;
  assign new_n8851_ = new_n8850_;
  assign new_n8852_ = new_n8851_;
  assign new_n8853_ = new_n8852_;
  assign new_n8854_ = new_n8851_;
  assign new_n8855_ = new_n8850_;
  assign new_n8856_ = new_n8855_;
  assign new_n8857_ = new_n8855_;
  assign new_n8858_ = new_n8833_;
  assign new_n8859_ = new_n8858_;
  assign new_n8860_ = new_n8859_;
  assign new_n8861_ = new_n8860_;
  assign new_n8862_ = new_n8860_;
  assign new_n8863_ = new_n8859_;
  assign new_n8864_ = new_n8863_;
  assign new_n8865_ = new_n8863_;
  assign new_n8866_ = new_n8858_;
  assign new_n8867_ = new_n8866_;
  assign new_n8868_ = new_n8867_;
  assign new_n8869_ = new_n8867_;
  assign new_n8870_ = new_n8866_;
  assign new_n8871_ = new_n8870_;
  assign new_n8872_ = new_n8870_;
  assign new_n8873_ = new_n3814_;
  assign new_n8874_ = new_n8873_;
  assign new_n8875_ = new_n8874_;
  assign new_n8876_ = new_n8875_;
  assign new_n8877_ = new_n8876_;
  assign new_n8878_ = new_n8877_;
  assign new_n8879_ = new_n8877_;
  assign new_n8880_ = new_n8876_;
  assign new_n8881_ = new_n8880_;
  assign new_n8882_ = new_n8880_;
  assign new_n8883_ = new_n8875_;
  assign new_n8884_ = new_n8883_;
  assign new_n8885_ = new_n8884_;
  assign new_n8886_ = new_n8884_;
  assign new_n8887_ = new_n8883_;
  assign new_n8888_ = new_n8887_;
  assign new_n8889_ = new_n8887_;
  assign new_n8890_ = new_n8874_;
  assign new_n8891_ = new_n8890_;
  assign new_n8892_ = new_n8891_;
  assign new_n8893_ = new_n8892_;
  assign new_n8894_ = new_n8891_;
  assign new_n8895_ = new_n8890_;
  assign new_n8896_ = new_n8895_;
  assign new_n8897_ = new_n8895_;
  assign new_n8898_ = new_n8873_;
  assign new_n8899_ = new_n8898_;
  assign new_n8900_ = new_n8899_;
  assign new_n8901_ = new_n8900_;
  assign new_n8902_ = new_n8900_;
  assign new_n8903_ = new_n8899_;
  assign new_n8904_ = new_n8903_;
  assign new_n8905_ = new_n8903_;
  assign new_n8906_ = new_n8898_;
  assign new_n8907_ = new_n8906_;
  assign new_n8908_ = new_n8907_;
  assign new_n8909_ = new_n8907_;
  assign new_n8910_ = new_n8906_;
  assign new_n8911_ = new_n8910_;
  assign new_n8912_ = new_n8910_;
  assign new_n8913_ = new_n2850_;
  assign new_n8914_ = new_n8913_;
  assign new_n8915_ = new_n2851_;
  assign new_n8916_ = new_n8915_;
  assign new_n8917_ = new_n5161_;
  assign new_n8918_ = new_n3807_;
  assign new_n8919_ = new_n8918_;
  assign new_n8920_ = new_n8919_;
  assign new_n8921_ = new_n8920_;
  assign new_n8922_ = new_n8921_;
  assign new_n8923_ = new_n8921_;
  assign new_n8924_ = new_n8920_;
  assign new_n8925_ = new_n8924_;
  assign new_n8926_ = new_n8924_;
  assign new_n8927_ = new_n8919_;
  assign new_n8928_ = new_n8927_;
  assign new_n8929_ = new_n8928_;
  assign new_n8930_ = new_n8928_;
  assign new_n8931_ = new_n8927_;
  assign new_n8932_ = new_n8931_;
  assign new_n8933_ = new_n8931_;
  assign new_n8934_ = new_n8918_;
  assign new_n8935_ = new_n8934_;
  assign new_n8936_ = new_n8935_;
  assign new_n8937_ = new_n8935_;
  assign new_n8938_ = new_n8934_;
  assign new_n8939_ = new_n8938_;
  assign new_n8940_ = new_n8938_;
  assign new_n8941_ = new_n3815_;
  assign new_n8942_ = new_n8941_;
  assign new_n8943_ = new_n8942_;
  assign new_n8944_ = new_n8943_;
  assign new_n8945_ = new_n8944_;
  assign new_n8946_ = new_n8944_;
  assign new_n8947_ = new_n8943_;
  assign new_n8948_ = new_n8947_;
  assign new_n8949_ = new_n8947_;
  assign new_n8950_ = new_n8942_;
  assign new_n8951_ = new_n8950_;
  assign new_n8952_ = new_n8951_;
  assign new_n8953_ = new_n8951_;
  assign new_n8954_ = new_n8950_;
  assign new_n8955_ = new_n8954_;
  assign new_n8956_ = new_n8954_;
  assign new_n8957_ = new_n8941_;
  assign new_n8958_ = new_n8957_;
  assign new_n8959_ = new_n8958_;
  assign new_n8960_ = new_n8958_;
  assign new_n8961_ = new_n8957_;
  assign new_n8962_ = new_n8961_;
  assign new_n8963_ = new_n8961_;
  assign new_n8964_ = new_n5171_;
  assign new_n8965_ = new_n8964_;
  assign new_n8966_ = new_n5170_;
  assign new_n8967_ = new_n8966_;
  assign new_n8968_ = new_n5176_;
  assign new_n8969_ = new_n2698_;
  assign new_n8970_ = new_n8969_;
  assign new_n8971_ = new_n2699_;
  assign new_n8972_ = new_n8971_;
  assign new_n8973_ = new_n5187_;
  assign new_n8974_ = new_n4404_;
  assign new_n8975_ = new_n4399_;
  assign new_n8976_ = new_n4405_;
  assign new_n8977_ = new_n4398_;
  assign new_n8978_ = new_n5202_;
  assign new_n8979_ = new_n8978_;
  assign new_n8980_ = new_n8979_;
  assign new_n8981_ = new_n8978_;
  assign new_n8982_ = new_n5203_;
  assign new_n8983_ = new_n8982_;
  assign new_n8984_ = new_n8983_;
  assign new_n8985_ = new_n8982_;
  assign new_n8986_ = new_n5210_;
  assign new_n8987_ = new_n5211_;
  assign new_n8988_ = new_n4211_;
  assign new_n8989_ = new_n5167_;
  assign new_n8990_ = new_n8989_;
  assign new_n8991_ = new_n8990_;
  assign new_n8992_ = new_n8989_;
  assign new_n8993_ = new_n3782_;
  assign new_n8994_ = new_n8993_;
  assign new_n8995_ = new_n8994_;
  assign new_n8996_ = new_n8995_;
  assign new_n8997_ = new_n8996_;
  assign new_n8998_ = new_n8996_;
  assign new_n8999_ = new_n8995_;
  assign new_n9000_ = new_n8999_;
  assign new_n9001_ = new_n8999_;
  assign new_n9002_ = new_n8994_;
  assign new_n9003_ = new_n9002_;
  assign new_n9004_ = new_n9002_;
  assign new_n9005_ = new_n8993_;
  assign new_n9006_ = new_n9005_;
  assign new_n9007_ = new_n9006_;
  assign new_n9008_ = new_n9006_;
  assign new_n9009_ = new_n9005_;
  assign new_n9010_ = new_n9009_;
  assign new_n9011_ = new_n9009_;
  assign new_n9012_ = new_n3774_;
  assign new_n9013_ = new_n9012_;
  assign new_n9014_ = new_n9013_;
  assign new_n9015_ = new_n9014_;
  assign new_n9016_ = new_n9015_;
  assign new_n9017_ = new_n9015_;
  assign new_n9018_ = new_n9014_;
  assign new_n9019_ = new_n9018_;
  assign new_n9020_ = new_n9018_;
  assign new_n9021_ = new_n9013_;
  assign new_n9022_ = new_n9021_;
  assign new_n9023_ = new_n9021_;
  assign new_n9024_ = new_n9012_;
  assign new_n9025_ = new_n9024_;
  assign new_n9026_ = new_n9025_;
  assign new_n9027_ = new_n9025_;
  assign new_n9028_ = new_n9024_;
  assign new_n9029_ = new_n9028_;
  assign new_n9030_ = new_n9028_;
  assign new_n9031_ = new_n5193_;
  assign new_n9032_ = new_n9031_;
  assign new_n9033_ = new_n9032_;
  assign new_n9034_ = new_n9031_;
  assign new_n9035_ = new_n3783_;
  assign new_n9036_ = new_n9035_;
  assign new_n9037_ = new_n9036_;
  assign new_n9038_ = new_n9037_;
  assign new_n9039_ = new_n9038_;
  assign new_n9040_ = new_n9038_;
  assign new_n9041_ = new_n9037_;
  assign new_n9042_ = new_n9041_;
  assign new_n9043_ = new_n9041_;
  assign new_n9044_ = new_n9036_;
  assign new_n9045_ = new_n9044_;
  assign new_n9046_ = new_n9044_;
  assign new_n9047_ = new_n9035_;
  assign new_n9048_ = new_n9047_;
  assign new_n9049_ = new_n9048_;
  assign new_n9050_ = new_n9048_;
  assign new_n9051_ = new_n9047_;
  assign new_n9052_ = new_n9051_;
  assign new_n9053_ = new_n9051_;
  assign new_n9054_ = new_n2706_;
  assign new_n9055_ = new_n3775_;
  assign new_n9056_ = new_n9055_;
  assign new_n9057_ = new_n9056_;
  assign new_n9058_ = new_n9057_;
  assign new_n9059_ = new_n9058_;
  assign new_n9060_ = new_n9058_;
  assign new_n9061_ = new_n9057_;
  assign new_n9062_ = new_n9061_;
  assign new_n9063_ = new_n9061_;
  assign new_n9064_ = new_n9056_;
  assign new_n9065_ = new_n9064_;
  assign new_n9066_ = new_n9064_;
  assign new_n9067_ = new_n9055_;
  assign new_n9068_ = new_n9067_;
  assign new_n9069_ = new_n9068_;
  assign new_n9070_ = new_n9068_;
  assign new_n9071_ = new_n9067_;
  assign new_n9072_ = new_n9071_;
  assign new_n9073_ = new_n9071_;
  assign new_n9074_ = new_n2858_;
  assign new_n9075_ = new_n5237_;
  assign new_n9076_ = new_n5238_;
  assign new_n9077_ = new_n5241_;
  assign new_n9078_ = new_n5242_;
  assign new_n9079_ = new_n5247_;
  assign new_n9080_ = new_n5248_;
  assign new_n9081_ = new_n5261_;
  assign new_n9082_ = new_n5278_;
  assign new_n9083_ = new_n5297_;
  assign new_n9084_ = new_n3790_;
  assign new_n9085_ = new_n9084_;
  assign new_n9086_ = new_n9085_;
  assign new_n9087_ = new_n9086_;
  assign new_n9088_ = new_n9087_;
  assign new_n9089_ = new_n9087_;
  assign new_n9090_ = new_n9086_;
  assign new_n9091_ = new_n9090_;
  assign new_n9092_ = new_n9090_;
  assign new_n9093_ = new_n9085_;
  assign new_n9094_ = new_n9093_;
  assign new_n9095_ = new_n9093_;
  assign new_n9096_ = new_n9084_;
  assign new_n9097_ = new_n9096_;
  assign new_n9098_ = new_n9097_;
  assign new_n9099_ = new_n9097_;
  assign new_n9100_ = new_n9096_;
  assign new_n9101_ = new_n9100_;
  assign new_n9102_ = new_n9100_;
  assign new_n9103_ = new_n3798_;
  assign new_n9104_ = new_n9103_;
  assign new_n9105_ = new_n9104_;
  assign new_n9106_ = new_n9105_;
  assign new_n9107_ = new_n9106_;
  assign new_n9108_ = new_n9106_;
  assign new_n9109_ = new_n9105_;
  assign new_n9110_ = new_n9109_;
  assign new_n9111_ = new_n9109_;
  assign new_n9112_ = new_n9104_;
  assign new_n9113_ = new_n9112_;
  assign new_n9114_ = new_n9112_;
  assign new_n9115_ = new_n9103_;
  assign new_n9116_ = new_n9115_;
  assign new_n9117_ = new_n9116_;
  assign new_n9118_ = new_n9116_;
  assign new_n9119_ = new_n9115_;
  assign new_n9120_ = new_n9119_;
  assign new_n9121_ = new_n9119_;
  assign new_n9122_ = new_n3791_;
  assign new_n9123_ = new_n9122_;
  assign new_n9124_ = new_n9123_;
  assign new_n9125_ = new_n9124_;
  assign new_n9126_ = new_n9125_;
  assign new_n9127_ = new_n9125_;
  assign new_n9128_ = new_n9124_;
  assign new_n9129_ = new_n9128_;
  assign new_n9130_ = new_n9128_;
  assign new_n9131_ = new_n9123_;
  assign new_n9132_ = new_n9131_;
  assign new_n9133_ = new_n9131_;
  assign new_n9134_ = new_n9122_;
  assign new_n9135_ = new_n9134_;
  assign new_n9136_ = new_n9135_;
  assign new_n9137_ = new_n9135_;
  assign new_n9138_ = new_n9134_;
  assign new_n9139_ = new_n9138_;
  assign new_n9140_ = new_n9138_;
  assign new_n9141_ = new_n3799_;
  assign new_n9142_ = new_n9141_;
  assign new_n9143_ = new_n9142_;
  assign new_n9144_ = new_n9143_;
  assign new_n9145_ = new_n9144_;
  assign new_n9146_ = new_n9144_;
  assign new_n9147_ = new_n9143_;
  assign new_n9148_ = new_n9147_;
  assign new_n9149_ = new_n9147_;
  assign new_n9150_ = new_n9142_;
  assign new_n9151_ = new_n9150_;
  assign new_n9152_ = new_n9150_;
  assign new_n9153_ = new_n9141_;
  assign new_n9154_ = new_n9153_;
  assign new_n9155_ = new_n9154_;
  assign new_n9156_ = new_n9154_;
  assign new_n9157_ = new_n9153_;
  assign new_n9158_ = new_n9157_;
  assign new_n9159_ = new_n9157_;
  assign new_n9160_ = new_n5319_;
  assign new_n9161_ = new_n5320_;
  assign new_n9162_ = new_n5323_;
  assign new_n9163_ = new_n5324_;
  assign new_n9164_ = new_n5327_;
  assign new_n9165_ = new_n9164_;
  assign new_n9166_ = new_n5328_;
  assign new_n9167_ = new_n9166_;
  assign new_n9168_ = new_n5331_;
  assign new_n9169_ = new_n5332_;
  assign new_n9170_ = new_n5345_;
  assign new_n9171_ = new_n5362_;
  assign new_n9172_ = new_n5381_;
  assign new_n9173_ = new_n5394_;
  assign new_n9174_ = new_n5411_;
  assign new_n9175_ = new_n5406_;
  assign new_n9176_ = new_n5412_;
  assign new_n9177_ = new_n5405_;
  assign new_n9178_ = new_n5421_;
  assign new_n9179_ = new_n9178_;
  assign new_n9180_ = new_n9178_;
  assign new_n9181_ = new_n5420_;
  assign new_n9182_ = new_n9181_;
  assign new_n9183_ = new_n9181_;
  assign new_n9184_ = new_n5422_;
  assign new_n9185_ = new_n9184_;
  assign new_n9186_ = new_n9184_;
  assign new_n9187_ = new_n5419_;
  assign new_n9188_ = new_n9187_;
  assign new_n9189_ = new_n9187_;
  assign new_n9190_ = new_n4428_;
  assign new_n9191_ = new_n9190_;
  assign new_n9192_ = new_n9190_;
  assign new_n9193_ = new_n4429_;
  assign new_n9194_ = new_n9193_;
  assign new_n9195_ = new_n9193_;
  assign new_n9196_ = new_n5458_;
  assign new_n9197_ = new_n5453_;
  assign new_n9198_ = new_n5459_;
  assign new_n9199_ = new_n5452_;
  assign new_n9200_ = new_n5468_;
  assign new_n9201_ = new_n9200_;
  assign new_n9202_ = new_n9200_;
  assign new_n9203_ = new_n5467_;
  assign new_n9204_ = new_n9203_;
  assign new_n9205_ = new_n9203_;
  assign new_n9206_ = new_n5469_;
  assign new_n9207_ = new_n9206_;
  assign new_n9208_ = new_n9206_;
  assign new_n9209_ = new_n5466_;
  assign new_n9210_ = new_n9209_;
  assign new_n9211_ = new_n9209_;
  assign new_n9212_ = new_n4431_;
  assign new_n9213_ = new_n9212_;
  assign new_n9214_ = new_n9212_;
  assign new_n9215_ = new_n4430_;
  assign new_n9216_ = new_n9215_;
  assign new_n9217_ = new_n9215_;
  assign new_n9218_ = new_n5497_;
  assign new_n9219_ = new_n9218_;
  assign new_n9220_ = new_n9218_;
  assign new_n9221_ = new_n5498_;
  assign new_n9222_ = new_n9221_;
  assign new_n9223_ = new_n9221_;
  assign new_n9224_ = new_n5501_;
  assign new_n9225_ = new_n5510_;
  assign new_n9226_ = new_n5523_;
  assign new_n9227_ = new_n5538_;
  assign new_n9228_ = new_n5549_;
  assign new_n9229_ = new_n5558_;
  assign new_n9230_ = new_n5571_;
  assign new_n9231_ = new_n5221_;
  assign new_n9232_ = new_n9231_;
  assign new_n9233_ = new_n9231_;
  assign new_n9234_ = new_n3664_;
  assign new_n9235_ = new_n9234_;
  assign new_n9236_ = new_n9235_;
  assign new_n9237_ = new_n9236_;
  assign new_n9238_ = new_n9237_;
  assign new_n9239_ = new_n9237_;
  assign new_n9240_ = new_n9236_;
  assign new_n9241_ = new_n9240_;
  assign new_n9242_ = new_n9240_;
  assign new_n9243_ = new_n9235_;
  assign new_n9244_ = new_n9243_;
  assign new_n9245_ = new_n9243_;
  assign new_n9246_ = new_n9234_;
  assign new_n9247_ = new_n9246_;
  assign new_n9248_ = new_n9247_;
  assign new_n9249_ = new_n9247_;
  assign new_n9250_ = new_n9246_;
  assign new_n9251_ = new_n9250_;
  assign new_n9252_ = new_n9250_;
  assign new_n9253_ = new_n3672_;
  assign new_n9254_ = new_n9253_;
  assign new_n9255_ = new_n9254_;
  assign new_n9256_ = new_n9255_;
  assign new_n9257_ = new_n9256_;
  assign new_n9258_ = new_n9256_;
  assign new_n9259_ = new_n9255_;
  assign new_n9260_ = new_n9259_;
  assign new_n9261_ = new_n9259_;
  assign new_n9262_ = new_n9254_;
  assign new_n9263_ = new_n9262_;
  assign new_n9264_ = new_n9262_;
  assign new_n9265_ = new_n9253_;
  assign new_n9266_ = new_n9265_;
  assign new_n9267_ = new_n9266_;
  assign new_n9268_ = new_n9266_;
  assign new_n9269_ = new_n9265_;
  assign new_n9270_ = new_n9269_;
  assign new_n9271_ = new_n9269_;
  assign new_n9272_ = new_n3665_;
  assign new_n9273_ = new_n9272_;
  assign new_n9274_ = new_n9273_;
  assign new_n9275_ = new_n9274_;
  assign new_n9276_ = new_n9275_;
  assign new_n9277_ = new_n9275_;
  assign new_n9278_ = new_n9274_;
  assign new_n9279_ = new_n9278_;
  assign new_n9280_ = new_n9278_;
  assign new_n9281_ = new_n9273_;
  assign new_n9282_ = new_n9281_;
  assign new_n9283_ = new_n9281_;
  assign new_n9284_ = new_n9272_;
  assign new_n9285_ = new_n9284_;
  assign new_n9286_ = new_n9285_;
  assign new_n9287_ = new_n9285_;
  assign new_n9288_ = new_n9284_;
  assign new_n9289_ = new_n9288_;
  assign new_n9290_ = new_n9288_;
  assign new_n9291_ = new_n3322_;
  assign new_n9292_ = new_n3673_;
  assign new_n9293_ = new_n9292_;
  assign new_n9294_ = new_n9293_;
  assign new_n9295_ = new_n9294_;
  assign new_n9296_ = new_n9295_;
  assign new_n9297_ = new_n9295_;
  assign new_n9298_ = new_n9294_;
  assign new_n9299_ = new_n9298_;
  assign new_n9300_ = new_n9298_;
  assign new_n9301_ = new_n9293_;
  assign new_n9302_ = new_n9301_;
  assign new_n9303_ = new_n9301_;
  assign new_n9304_ = new_n9292_;
  assign new_n9305_ = new_n9304_;
  assign new_n9306_ = new_n9305_;
  assign new_n9307_ = new_n9305_;
  assign new_n9308_ = new_n9304_;
  assign new_n9309_ = new_n9308_;
  assign new_n9310_ = new_n9308_;
  assign new_n9311_ = new_n3330_;
  assign new_n9312_ = new_n3194_;
  assign new_n9313_ = new_n9312_;
  assign new_n9314_ = new_n9313_;
  assign new_n9315_ = new_n9314_;
  assign new_n9316_ = new_n9315_;
  assign new_n9317_ = new_n9315_;
  assign new_n9318_ = new_n9314_;
  assign new_n9319_ = new_n9318_;
  assign new_n9320_ = new_n9318_;
  assign new_n9321_ = new_n9313_;
  assign new_n9322_ = new_n9321_;
  assign new_n9323_ = new_n9322_;
  assign new_n9324_ = new_n9321_;
  assign new_n9325_ = new_n9312_;
  assign new_n9326_ = new_n9325_;
  assign new_n9327_ = new_n9326_;
  assign new_n9328_ = new_n9326_;
  assign new_n9329_ = new_n9325_;
  assign new_n9330_ = new_n9329_;
  assign new_n9331_ = new_n9329_;
  assign new_n9332_ = new_n3680_;
  assign new_n9333_ = new_n9332_;
  assign new_n9334_ = new_n9333_;
  assign new_n9335_ = new_n9334_;
  assign new_n9336_ = new_n9335_;
  assign new_n9337_ = new_n9335_;
  assign new_n9338_ = new_n9334_;
  assign new_n9339_ = new_n9338_;
  assign new_n9340_ = new_n9338_;
  assign new_n9341_ = new_n9333_;
  assign new_n9342_ = new_n9341_;
  assign new_n9343_ = new_n9341_;
  assign new_n9344_ = new_n9332_;
  assign new_n9345_ = new_n9344_;
  assign new_n9346_ = new_n9345_;
  assign new_n9347_ = new_n9345_;
  assign new_n9348_ = new_n9344_;
  assign new_n9349_ = new_n9348_;
  assign new_n9350_ = new_n9348_;
  assign new_n9351_ = new_n3688_;
  assign new_n9352_ = new_n9351_;
  assign new_n9353_ = new_n9352_;
  assign new_n9354_ = new_n9353_;
  assign new_n9355_ = new_n9354_;
  assign new_n9356_ = new_n9354_;
  assign new_n9357_ = new_n9353_;
  assign new_n9358_ = new_n9357_;
  assign new_n9359_ = new_n9357_;
  assign new_n9360_ = new_n9352_;
  assign new_n9361_ = new_n9360_;
  assign new_n9362_ = new_n9360_;
  assign new_n9363_ = new_n9351_;
  assign new_n9364_ = new_n9363_;
  assign new_n9365_ = new_n9364_;
  assign new_n9366_ = new_n9364_;
  assign new_n9367_ = new_n9363_;
  assign new_n9368_ = new_n9367_;
  assign new_n9369_ = new_n9367_;
  assign new_n9370_ = new_n3681_;
  assign new_n9371_ = new_n9370_;
  assign new_n9372_ = new_n9371_;
  assign new_n9373_ = new_n9372_;
  assign new_n9374_ = new_n9373_;
  assign new_n9375_ = new_n9373_;
  assign new_n9376_ = new_n9372_;
  assign new_n9377_ = new_n9376_;
  assign new_n9378_ = new_n9376_;
  assign new_n9379_ = new_n9371_;
  assign new_n9380_ = new_n9379_;
  assign new_n9381_ = new_n9379_;
  assign new_n9382_ = new_n9370_;
  assign new_n9383_ = new_n9382_;
  assign new_n9384_ = new_n9383_;
  assign new_n9385_ = new_n9383_;
  assign new_n9386_ = new_n9382_;
  assign new_n9387_ = new_n9386_;
  assign new_n9388_ = new_n9386_;
  assign new_n9389_ = new_n3689_;
  assign new_n9390_ = new_n9389_;
  assign new_n9391_ = new_n9390_;
  assign new_n9392_ = new_n9391_;
  assign new_n9393_ = new_n9392_;
  assign new_n9394_ = new_n9392_;
  assign new_n9395_ = new_n9391_;
  assign new_n9396_ = new_n9395_;
  assign new_n9397_ = new_n9395_;
  assign new_n9398_ = new_n9390_;
  assign new_n9399_ = new_n9398_;
  assign new_n9400_ = new_n9398_;
  assign new_n9401_ = new_n9389_;
  assign new_n9402_ = new_n9401_;
  assign new_n9403_ = new_n9402_;
  assign new_n9404_ = new_n9402_;
  assign new_n9405_ = new_n9401_;
  assign new_n9406_ = new_n9405_;
  assign new_n9407_ = new_n9405_;
  assign new_n9408_ = new_n5267_;
  assign new_n9409_ = new_n9408_;
  assign new_n9410_ = new_n9409_;
  assign new_n9411_ = new_n9408_;
  assign new_n9412_ = new_n5351_;
  assign new_n9413_ = new_n9412_;
  assign new_n9414_ = new_n9413_;
  assign new_n9415_ = new_n9412_;
  assign new_n9416_ = new_n2810_;
  assign new_n9417_ = new_n2794_;
  assign new_n9418_ = new_n5284_;
  assign new_n9419_ = new_n9418_;
  assign new_n9420_ = new_n9419_;
  assign new_n9421_ = new_n9418_;
  assign new_n9422_ = new_n5368_;
  assign new_n9423_ = new_n9422_;
  assign new_n9424_ = new_n9423_;
  assign new_n9425_ = new_n9422_;
  assign new_n9426_ = new_n2898_;
  assign new_n9427_ = new_n2730_;
  assign new_n9428_ = new_n5303_;
  assign new_n9429_ = new_n9428_;
  assign new_n9430_ = new_n9429_;
  assign new_n9431_ = new_n9428_;
  assign new_n9432_ = new_n5387_;
  assign new_n9433_ = new_n9432_;
  assign new_n9434_ = new_n9433_;
  assign new_n9435_ = new_n9432_;
  assign new_n9436_ = new_n2890_;
  assign new_n9437_ = new_n2722_;
  assign new_n9438_ = new_n5182_;
  assign new_n9439_ = new_n9438_;
  assign new_n9440_ = new_n9439_;
  assign new_n9441_ = new_n9438_;
  assign new_n9442_ = new_n5400_;
  assign new_n9443_ = new_n9442_;
  assign new_n9444_ = new_n9443_;
  assign new_n9445_ = new_n9442_;
  assign new_n9446_ = new_n2874_;
  assign new_n9447_ = new_n2882_;
  assign new_n9448_ = new_n3370_;
  assign new_n9449_ = new_n3290_;
  assign new_n9450_ = new_n3338_;
  assign new_n9451_ = new_n3258_;
  assign new_n9452_ = new_n3250_;
  assign new_n9453_ = new_n3242_;
  assign new_n9454_ = new_n3234_;
  assign new_n9455_ = new_n3226_;
  assign new_n9456_ = new_n4792_;
  assign new_n9457_ = new_n3767_;
  assign new_n9458_ = new_n3759_;
  assign new_n9459_ = new_n3902_;
  assign new_n9460_ = new_n3170_;
  assign new_n9461_ = new_n3171_;
  assign new_n9462_ = new_n5792_;
  assign new_n9463_ = new_n5791_;
  assign new_n9464_ = new_n5798_;
  assign new_n9465_ = new_n3766_;
  assign new_n9466_ = new_n3114_;
  assign new_n9467_ = new_n3758_;
  assign new_n9468_ = new_n5220_;
  assign new_n9469_ = new_n5809_;
  assign new_n9470_ = new_n3643_;
  assign new_n9471_ = new_n3627_;
  assign new_n9472_ = new_n5447_;
  assign new_n9473_ = new_n3651_;
  assign new_n9474_ = new_n5494_;
  assign new_n9475_ = new_n5001_;
  assign new_n9476_ = new_n5048_;
  assign new_n9477_ = new_n3427_;
  assign new_n9478_ = new_n3855_;
  assign new_n9479_ = new_n3854_;
  assign new_n9480_ = new_n5820_;
  assign new_n9481_ = new_n9480_;
  assign new_n9482_ = new_n9481_;
  assign new_n9483_ = new_n9480_;
  assign new_n9484_ = new_n5871_;
  assign new_n9485_ = new_n9484_;
  assign new_n9486_ = new_n9485_;
  assign new_n9487_ = new_n9484_;
  assign new_n9488_ = new_n3018_;
  assign new_n9489_ = new_n3010_;
  assign new_n9490_ = new_n5828_;
  assign new_n9491_ = new_n9490_;
  assign new_n9492_ = new_n9491_;
  assign new_n9493_ = new_n9490_;
  assign new_n9494_ = new_n5879_;
  assign new_n9495_ = new_n9494_;
  assign new_n9496_ = new_n9495_;
  assign new_n9497_ = new_n9494_;
  assign new_n9498_ = new_n2818_;
  assign new_n9499_ = new_n2826_;
  assign new_n9500_ = new_n5836_;
  assign new_n9501_ = new_n9500_;
  assign new_n9502_ = new_n9501_;
  assign new_n9503_ = new_n9500_;
  assign new_n9504_ = new_n5887_;
  assign new_n9505_ = new_n9504_;
  assign new_n9506_ = new_n9505_;
  assign new_n9507_ = new_n9504_;
  assign new_n9508_ = new_n2994_;
  assign new_n9509_ = new_n3002_;
  assign new_n9510_ = new_n5844_;
  assign new_n9511_ = new_n9510_;
  assign new_n9512_ = new_n9511_;
  assign new_n9513_ = new_n9510_;
  assign new_n9514_ = new_n5895_;
  assign new_n9515_ = new_n9514_;
  assign new_n9516_ = new_n9515_;
  assign new_n9517_ = new_n9514_;
  assign new_n9518_ = new_n2970_;
  assign new_n9519_ = new_n2802_;
  assign new_n9520_ = new_n3378_;
  assign new_n9521_ = new_n3298_;
  assign new_n9522_ = new_n3362_;
  assign new_n9523_ = new_n3282_;
  assign new_n9524_ = new_n3354_;
  assign new_n9525_ = new_n3274_;
  assign new_n9526_ = new_n3346_;
  assign new_n9527_ = new_n3266_;
  assign new_n9528_ = new_n6082_;
  assign new_n9529_ = new_n6087_;
  assign new_n9530_ = new_n6092_;
  assign new_n9531_ = new_n6098_;
  assign new_n9532_ = new_n6103_;
  assign new_n9533_ = new_n6116_;
  assign new_n9534_ = new_n9533_;
  assign new_n9535_ = new_n9533_;
  assign new_n9536_ = new_n6124_;
  assign new_n9537_ = new_n9536_;
  assign new_n9538_ = new_n9536_;
  assign new_n9539_ = new_n2714_;
  assign new_n9540_ = new_n2866_;
  assign new_n9541_ = new_n3306_;
  assign new_n9542_ = new_n3314_;
  assign new_n9543_ = new_n4461_;
  assign new_n9544_ = new_n9543_;
  assign new_n9545_ = new_n9544_;
  assign new_n9546_ = new_n9544_;
  assign new_n9547_ = new_n9543_;
  assign new_n9548_ = new_n9547_;
  assign new_n9549_ = new_n9547_;
  assign new_n9550_ = new_n4188_;
  assign new_n9551_ = new_n9550_;
  assign new_n9552_ = new_n9551_;
  assign new_n9553_ = new_n9550_;
  assign new_n9554_ = new_n4460_;
  assign new_n9555_ = new_n9554_;
  assign new_n9556_ = new_n9555_;
  assign new_n9557_ = new_n9556_;
  assign new_n9558_ = new_n9555_;
  assign new_n9559_ = new_n9554_;
  assign new_n9560_ = new_n9559_;
  assign new_n9561_ = new_n9559_;
  assign new_n9562_ = new_n4189_;
  assign new_n9563_ = new_n9562_;
  assign new_n9564_ = new_n9562_;
  assign new_n9565_ = new_n4465_;
  assign new_n9566_ = new_n9565_;
  assign new_n9567_ = new_n9566_;
  assign new_n9568_ = new_n9566_;
  assign new_n9569_ = new_n9565_;
  assign new_n9570_ = new_n9569_;
  assign new_n9571_ = new_n4464_;
  assign new_n9572_ = new_n9571_;
  assign new_n9573_ = new_n9572_;
  assign new_n9574_ = new_n9572_;
  assign new_n9575_ = new_n9571_;
  assign new_n9576_ = new_n9575_;
  assign new_n9577_ = new_n9575_;
  assign new_n9578_ = new_n4563_;
  assign new_n9579_ = new_n9578_;
  assign new_n9580_ = new_n9579_;
  assign new_n9581_ = new_n9579_;
  assign new_n9582_ = new_n9578_;
  assign new_n9583_ = new_n9582_;
  assign new_n9584_ = new_n9582_;
  assign new_n9585_ = new_n4546_;
  assign new_n9586_ = new_n4562_;
  assign new_n9587_ = new_n9586_;
  assign new_n9588_ = new_n9587_;
  assign new_n9589_ = new_n9588_;
  assign new_n9590_ = new_n9587_;
  assign new_n9591_ = new_n9586_;
  assign new_n9592_ = new_n9591_;
  assign new_n9593_ = new_n9591_;
  assign new_n9594_ = new_n4547_;
  assign new_n9595_ = new_n4565_;
  assign new_n9596_ = new_n9595_;
  assign new_n9597_ = new_n9596_;
  assign new_n9598_ = new_n9596_;
  assign new_n9599_ = new_n9595_;
  assign new_n9600_ = new_n9599_;
  assign new_n9601_ = new_n4564_;
  assign new_n9602_ = new_n9601_;
  assign new_n9603_ = new_n9602_;
  assign new_n9604_ = new_n9602_;
  assign new_n9605_ = new_n9601_;
  assign new_n9606_ = new_n9605_;
  assign new_n9607_ = new_n9605_;
  assign new_n9608_ = new_n3942_;
  assign new_n9609_ = new_n3943_;
  assign new_n9610_ = new_n3940_;
  assign new_n9611_ = new_n9610_;
  assign new_n9612_ = new_n9611_;
  assign new_n9613_ = new_n9611_;
  assign new_n9614_ = new_n9610_;
  assign new_n9615_ = new_n9614_;
  assign new_n9616_ = new_n3941_;
  assign new_n9617_ = new_n9616_;
  assign new_n9618_ = new_n9617_;
  assign new_n9619_ = new_n9617_;
  assign new_n9620_ = new_n9616_;
  assign new_n9621_ = new_n9620_;
  assign new_n9622_ = new_n4006_;
  assign new_n9623_ = new_n9622_;
  assign new_n9624_ = new_n9623_;
  assign new_n9625_ = new_n9623_;
  assign new_n9626_ = new_n9622_;
  assign new_n9627_ = new_n4007_;
  assign new_n9628_ = new_n9627_;
  assign new_n9629_ = new_n9628_;
  assign new_n9630_ = new_n9628_;
  assign new_n9631_ = new_n9627_;
  assign new_n9632_ = new_n4230_;
  assign new_n9633_ = new_n9632_;
  assign new_n9634_ = new_n9633_;
  assign new_n9635_ = new_n9632_;
  assign new_n9636_ = new_n4231_;
  assign new_n9637_ = new_n9636_;
  assign new_n9638_ = new_n9637_;
  assign new_n9639_ = new_n9636_;
  assign new_n9640_ = new_n3946_;
  assign new_n9641_ = new_n3947_;
  assign new_n9642_ = new_n3944_;
  assign new_n9643_ = new_n9642_;
  assign new_n9644_ = new_n9643_;
  assign new_n9645_ = new_n9643_;
  assign new_n9646_ = new_n9642_;
  assign new_n9647_ = new_n9646_;
  assign new_n9648_ = new_n3945_;
  assign new_n9649_ = new_n9648_;
  assign new_n9650_ = new_n9649_;
  assign new_n9651_ = new_n9649_;
  assign new_n9652_ = new_n9648_;
  assign new_n9653_ = new_n9652_;
  assign new_n9654_ = new_n4012_;
  assign new_n9655_ = new_n9654_;
  assign new_n9656_ = new_n9655_;
  assign new_n9657_ = new_n9655_;
  assign new_n9658_ = new_n9654_;
  assign new_n9659_ = new_n4013_;
  assign new_n9660_ = new_n9659_;
  assign new_n9661_ = new_n9660_;
  assign new_n9662_ = new_n9660_;
  assign new_n9663_ = new_n9659_;
  assign new_n9664_ = new_n4232_;
  assign new_n9665_ = new_n9664_;
  assign new_n9666_ = new_n9665_;
  assign new_n9667_ = new_n9664_;
  assign new_n9668_ = new_n4233_;
  assign new_n9669_ = new_n9668_;
  assign new_n9670_ = new_n9669_;
  assign new_n9671_ = new_n9668_;
  assign new_n9672_ = new_n4088_;
  assign new_n9673_ = new_n9672_;
  assign new_n9674_ = new_n9672_;
  assign new_n9675_ = new_n4082_;
  assign new_n9676_ = new_n9675_;
  assign new_n9677_ = new_n9675_;
  assign new_n9678_ = new_n4089_;
  assign new_n9679_ = new_n9678_;
  assign new_n9680_ = new_n4083_;
  assign new_n9681_ = new_n9680_;
  assign new_n9682_ = new_n4086_;
  assign new_n9683_ = new_n9682_;
  assign new_n9684_ = new_n9682_;
  assign new_n9685_ = new_n4084_;
  assign new_n9686_ = new_n9685_;
  assign new_n9687_ = new_n9685_;
  assign new_n9688_ = new_n4087_;
  assign new_n9689_ = new_n9688_;
  assign new_n9690_ = new_n4085_;
  assign new_n9691_ = new_n9690_;
  assign new_n9692_ = new_n3913_;
  assign new_n9693_ = new_n9692_;
  assign new_n9694_ = new_n3912_;
  assign new_n9695_ = new_n9694_;
  assign new_n9696_ = new_n9694_;
  assign new_n9697_ = new_n4482_;
  assign new_n9698_ = new_n4480_;
  assign new_n9699_ = new_n4134_;
  assign new_n9700_ = new_n3496_;
  assign new_n9701_ = new_n9700_;
  assign new_n9702_ = new_n9701_;
  assign new_n9703_ = new_n9700_;
  assign new_n9704_ = new_n3497_;
  assign new_n9705_ = new_n4099_;
  assign new_n9706_ = new_n4136_;
  assign new_n9707_ = new_n3408_;
  assign new_n9708_ = new_n9707_;
  assign new_n9709_ = new_n9708_;
  assign new_n9710_ = new_n9707_;
  assign new_n9711_ = new_n3409_;
  assign new_n9712_ = new_n4101_;
  assign new_n9713_ = new_n4688_;
  assign new_n9714_ = new_n4504_;
  assign new_n9715_ = new_n9714_;
  assign new_n9716_ = new_n4505_;
  assign new_n9717_ = new_n4690_;
  assign new_n9718_ = new_n4257_;
  assign new_n9719_ = new_n4256_;
  assign new_n9720_ = new_n9719_;
  assign new_n9721_ = new_n3982_;
  assign new_n9722_ = new_n9721_;
  assign new_n9723_ = new_n9721_;
  assign new_n9724_ = new_n3976_;
  assign new_n9725_ = new_n9724_;
  assign new_n9726_ = new_n9725_;
  assign new_n9727_ = new_n9725_;
  assign new_n9728_ = new_n9724_;
  assign new_n9729_ = new_n9728_;
  assign new_n9730_ = new_n3974_;
  assign new_n9731_ = new_n9730_;
  assign new_n9732_ = new_n3962_;
  assign new_n9733_ = new_n9732_;
  assign new_n9734_ = new_n9733_;
  assign new_n9735_ = new_n9733_;
  assign new_n9736_ = new_n9732_;
  assign new_n9737_ = new_n3973_;
  assign new_n9738_ = new_n9737_;
  assign new_n9739_ = new_n3965_;
  assign new_n9740_ = new_n9739_;
  assign new_n9741_ = new_n9740_;
  assign new_n9742_ = new_n9740_;
  assign new_n9743_ = new_n9739_;
  assign new_n9744_ = new_n3981_;
  assign new_n9745_ = new_n3979_;
  assign new_n9746_ = new_n9745_;
  assign new_n9747_ = new_n9746_;
  assign new_n9748_ = new_n9745_;
  assign new_n9749_ = new_n4676_;
  assign new_n9750_ = new_n4672_;
  assign new_n9751_ = new_n4680_;
  assign new_n9752_ = new_n4668_;
  assign new_n9753_ = new_n4004_;
  assign new_n9754_ = new_n9753_;
  assign new_n9755_ = new_n3991_;
  assign new_n9756_ = new_n9755_;
  assign new_n9757_ = new_n9755_;
  assign new_n9758_ = new_n4005_;
  assign new_n9759_ = new_n3990_;
  assign new_n9760_ = new_n9759_;
  assign new_n9761_ = new_n9760_;
  assign new_n9762_ = new_n9760_;
  assign new_n9763_ = new_n9759_;
  assign new_n9764_ = new_n3963_;
  assign new_n9765_ = new_n9764_;
  assign new_n9766_ = new_n9764_;
  assign new_n9767_ = new_n3975_;
  assign new_n9768_ = new_n3972_;
  assign new_n9769_ = new_n9768_;
  assign new_n9770_ = new_n9768_;
  assign new_n9771_ = new_n3964_;
  assign new_n9772_ = new_n9771_;
  assign new_n9773_ = new_n9772_;
  assign new_n9774_ = new_n9772_;
  assign new_n9775_ = new_n9771_;
  assign new_n9776_ = new_n4692_;
  assign new_n9777_ = new_n9776_;
  assign new_n9778_ = new_n9777_;
  assign new_n9779_ = new_n9776_;
  assign new_n9780_ = new_n4686_;
  assign new_n9781_ = new_n9780_;
  assign new_n9782_ = new_n9781_;
  assign new_n9783_ = new_n9780_;
  assign new_n9784_ = new_n4693_;
  assign new_n9785_ = new_n9784_;
  assign new_n9786_ = new_n9784_;
  assign new_n9787_ = new_n4687_;
  assign new_n9788_ = new_n9787_;
  assign new_n9789_ = new_n9787_;
  assign new_n9790_ = new_n4702_;
  assign new_n9791_ = new_n4699_;
  assign new_n9792_ = new_n4703_;
  assign new_n9793_ = new_n4698_;
  assign new_n9794_ = new_n4704_;
  assign new_n9795_ = new_n4701_;
  assign new_n9796_ = new_n4705_;
  assign new_n9797_ = new_n4700_;
  assign new_n9798_ = new_n4706_;
  assign new_n9799_ = new_n4695_;
  assign new_n9800_ = new_n4707_;
  assign new_n9801_ = new_n4694_;
  assign new_n9802_ = new_n4708_;
  assign new_n9803_ = new_n4697_;
  assign new_n9804_ = new_n4709_;
  assign new_n9805_ = new_n4696_;
  assign new_n9806_ = new_n4674_;
  assign new_n9807_ = new_n4670_;
  assign new_n9808_ = new_n4678_;
  assign new_n9809_ = new_n4666_;
  assign new_n9810_ = new_n3504_;
  assign new_n9811_ = new_n4506_;
  assign new_n9812_ = new_n3440_;
  assign new_n9813_ = new_n4258_;
  assign new_n9814_ = new_n4252_;
  assign new_n9815_ = new_n9814_;
  assign new_n9816_ = new_n9815_;
  assign new_n9817_ = new_n9815_;
  assign new_n9818_ = new_n9814_;
  assign new_n9819_ = new_n9818_;
  assign new_n9820_ = new_n3482_;
  assign new_n9821_ = new_n4253_;
  assign new_n9822_ = new_n9821_;
  assign new_n9823_ = new_n9822_;
  assign new_n9824_ = new_n9821_;
  assign new_n9825_ = new_n4254_;
  assign new_n9826_ = new_n9825_;
  assign new_n9827_ = new_n9826_;
  assign new_n9828_ = new_n9826_;
  assign new_n9829_ = new_n9825_;
  assign new_n9830_ = new_n9829_;
  assign new_n9831_ = new_n3394_;
  assign new_n9832_ = new_n4255_;
  assign new_n9833_ = new_n9832_;
  assign new_n9834_ = new_n9833_;
  assign new_n9835_ = new_n9832_;
  assign new_n9836_ = new_n6384_;
  assign new_n9837_ = new_n6169_;
  assign new_n9838_ = new_n9837_;
  assign new_n9839_ = new_n9837_;
  assign new_n9840_ = new_n6385_;
  assign new_n9841_ = new_n6170_;
  assign new_n9842_ = new_n9841_;
  assign new_n9843_ = new_n9842_;
  assign new_n9844_ = new_n9841_;
  assign new_n9845_ = new_n4040_;
  assign new_n9846_ = new_n9845_;
  assign new_n9847_ = new_n4041_;
  assign new_n9848_ = new_n6394_;
  assign new_n9849_ = new_n6236_;
  assign new_n9850_ = new_n9849_;
  assign new_n9851_ = new_n3656_;
  assign new_n9852_ = new_n9851_;
  assign new_n9853_ = new_n6401_;
  assign new_n9854_ = new_n6402_;
  assign new_n9855_ = new_n6411_;
  assign new_n9856_ = new_n6235_;
  assign new_n9857_ = new_n6197_;
  assign new_n9858_ = new_n3657_;
  assign new_n9859_ = new_n9858_;
  assign new_n9860_ = new_n6423_;
  assign new_n9861_ = new_n6424_;
  assign new_n9862_ = new_n6439_;
  assign new_n9863_ = new_n6440_;
  assign new_n9864_ = new_n6456_;
  assign new_n9865_ = new_n4578_;
  assign new_n9866_ = new_n9865_;
  assign new_n9867_ = new_n9866_;
  assign new_n9868_ = new_n9867_;
  assign new_n9869_ = new_n9867_;
  assign new_n9870_ = new_n9866_;
  assign new_n9871_ = new_n9865_;
  assign new_n9872_ = new_n9871_;
  assign new_n9873_ = new_n9871_;
  assign new_n9874_ = new_n6457_;
  assign new_n9875_ = new_n4579_;
  assign new_n9876_ = new_n9875_;
  assign new_n9877_ = new_n9875_;
  assign new_n9878_ = new_n4042_;
  assign new_n9879_ = new_n9878_;
  assign new_n9880_ = new_n4043_;
  assign new_n9881_ = new_n6466_;
  assign new_n9882_ = new_n6265_;
  assign new_n9883_ = new_n3695_;
  assign new_n9884_ = new_n9883_;
  assign new_n9885_ = new_n6473_;
  assign new_n9886_ = new_n6474_;
  assign new_n9887_ = new_n6483_;
  assign new_n9888_ = new_n6266_;
  assign new_n9889_ = new_n9888_;
  assign new_n9890_ = new_n6205_;
  assign new_n9891_ = new_n3694_;
  assign new_n9892_ = new_n9891_;
  assign new_n9893_ = new_n6495_;
  assign new_n9894_ = new_n6496_;
  assign new_n9895_ = new_n6511_;
  assign new_n9896_ = new_n6512_;
  assign new_n9897_ = new_n3977_;
  assign new_n9898_ = new_n9897_;
  assign new_n9899_ = new_n9897_;
  assign new_n9900_ = new_n3983_;
  assign new_n9901_ = new_n4228_;
  assign new_n9902_ = new_n9901_;
  assign new_n9903_ = new_n4229_;
  assign new_n9904_ = new_n3980_;
  assign new_n9905_ = new_n9904_;
  assign new_n9906_ = new_n9904_;
  assign new_n9907_ = new_n3978_;
  assign new_n9908_ = new_n9907_;
  assign new_n9909_ = new_n9908_;
  assign new_n9910_ = new_n9908_;
  assign new_n9911_ = new_n9907_;
  assign new_n9912_ = new_n3382_;
  assign new_n9913_ = new_n9912_;
  assign new_n9914_ = new_n9913_;
  assign new_n9915_ = new_n9912_;
  assign new_n9916_ = new_n3564_;
  assign new_n9917_ = new_n9916_;
  assign new_n9918_ = new_n9916_;
  assign new_n9919_ = new_n6294_;
  assign new_n9920_ = new_n3592_;
  assign new_n9921_ = new_n9920_;
  assign new_n9922_ = new_n9920_;
  assign new_n9923_ = new_n6288_;
  assign new_n9924_ = new_n3488_;
  assign new_n9925_ = new_n3400_;
  assign new_n9926_ = new_n3918_;
  assign new_n9927_ = new_n9926_;
  assign new_n9928_ = new_n9926_;
  assign new_n9929_ = new_n3916_;
  assign new_n9930_ = new_n9929_;
  assign new_n9931_ = new_n9930_;
  assign new_n9932_ = new_n9930_;
  assign new_n9933_ = new_n9929_;
  assign new_n9934_ = new_n3970_;
  assign new_n9935_ = new_n9934_;
  assign new_n9936_ = new_n9934_;
  assign new_n9937_ = new_n3960_;
  assign new_n9938_ = new_n9937_;
  assign new_n9939_ = new_n9937_;
  assign new_n9940_ = new_n3908_;
  assign new_n9941_ = new_n9940_;
  assign new_n9942_ = new_n9940_;
  assign new_n9943_ = new_n3894_;
  assign new_n9944_ = new_n9943_;
  assign new_n9945_ = new_n9944_;
  assign new_n9946_ = new_n9944_;
  assign new_n9947_ = new_n9943_;
  assign new_n9948_ = new_n3910_;
  assign new_n9949_ = new_n9948_;
  assign new_n9950_ = new_n9948_;
  assign new_n9951_ = new_n3896_;
  assign new_n9952_ = new_n9951_;
  assign new_n9953_ = new_n9952_;
  assign new_n9954_ = new_n9952_;
  assign new_n9955_ = new_n9951_;
  assign new_n9956_ = new_n3968_;
  assign new_n9957_ = new_n9956_;
  assign new_n9958_ = new_n3966_;
  assign new_n9959_ = new_n9958_;
  assign new_n9960_ = new_n9959_;
  assign new_n9961_ = new_n9958_;
  assign new_n9962_ = new_n3904_;
  assign new_n9963_ = new_n9962_;
  assign new_n9964_ = new_n3898_;
  assign new_n9965_ = new_n9964_;
  assign new_n9966_ = new_n9965_;
  assign new_n9967_ = new_n9965_;
  assign new_n9968_ = new_n9964_;
  assign new_n9969_ = new_n3906_;
  assign new_n9970_ = new_n9969_;
  assign new_n9971_ = new_n3900_;
  assign new_n9972_ = new_n9971_;
  assign new_n9973_ = new_n9972_;
  assign new_n9974_ = new_n9972_;
  assign new_n9975_ = new_n9971_;
  assign new_n9976_ = new_n3870_;
  assign new_n9977_ = new_n3868_;
  assign new_n9978_ = new_n3885_;
  assign new_n9979_ = new_n9978_;
  assign new_n9980_ = new_n9979_;
  assign new_n9981_ = new_n9978_;
  assign new_n9982_ = new_n3456_;
  assign new_n9983_ = new_n3884_;
  assign new_n9984_ = new_n9983_;
  assign new_n9985_ = new_n9984_;
  assign new_n9986_ = new_n9984_;
  assign new_n9987_ = new_n9983_;
  assign new_n9988_ = new_n3457_;
  assign new_n9989_ = new_n3876_;
  assign new_n9990_ = new_n3872_;
  assign new_n9991_ = new_n3524_;
  assign new_n9992_ = new_n6314_;
  assign new_n9993_ = new_n9992_;
  assign new_n9994_ = new_n9992_;
  assign new_n9995_ = new_n6301_;
  assign new_n9996_ = new_n6571_;
  assign new_n9997_ = new_n9996_;
  assign new_n9998_ = new_n6311_;
  assign new_n9999_ = new_n9998_;
  assign new_n10000_ = new_n9999_;
  assign new_n10001_ = new_n9998_;
  assign new_n10002_ = new_n6302_;
  assign new_n10003_ = new_n10002_;
  assign new_n10004_ = new_n6303_;
  assign new_n10005_ = new_n10004_;
  assign new_n10006_ = new_n4030_;
  assign new_n10007_ = new_n10006_;
  assign new_n10008_ = new_n10007_;
  assign new_n10009_ = new_n10007_;
  assign new_n10010_ = new_n10006_;
  assign new_n10011_ = new_n10010_;
  assign new_n10012_ = new_n10010_;
  assign new_n10013_ = new_n6304_;
  assign new_n10014_ = new_n6576_;
  assign new_n10015_ = new_n10014_;
  assign new_n10016_ = new_n3905_;
  assign new_n10017_ = new_n3907_;
  assign new_n10018_ = new_n6583_;
  assign new_n10019_ = new_n3924_;
  assign new_n10020_ = new_n10019_;
  assign new_n10021_ = new_n10019_;
  assign new_n10022_ = new_n6532_;
  assign new_n10023_ = new_n6320_;
  assign new_n10024_ = new_n10023_;
  assign new_n10025_ = new_n6588_;
  assign new_n10026_ = new_n6526_;
  assign new_n10027_ = new_n6592_;
  assign new_n10028_ = new_n6573_;
  assign new_n10029_ = new_n6379_;
  assign new_n10030_ = new_n6572_;
  assign new_n10031_ = new_n6575_;
  assign new_n10032_ = new_n6578_;
  assign new_n10033_ = new_n4036_;
  assign new_n10034_ = new_n3928_;
  assign new_n10035_ = new_n3917_;
  assign new_n10036_ = new_n10035_;
  assign new_n10037_ = new_n10035_;
  assign new_n10038_ = new_n3961_;
  assign new_n10039_ = new_n3895_;
  assign new_n10040_ = new_n10039_;
  assign new_n10041_ = new_n10039_;
  assign new_n10042_ = new_n3897_;
  assign new_n10043_ = new_n10042_;
  assign new_n10044_ = new_n10042_;
  assign new_n10045_ = new_n3967_;
  assign new_n10046_ = new_n10045_;
  assign new_n10047_ = new_n3969_;
  assign new_n10048_ = new_n3899_;
  assign new_n10049_ = new_n10048_;
  assign new_n10050_ = new_n10048_;
  assign new_n10051_ = new_n3901_;
  assign new_n10052_ = new_n10051_;
  assign new_n10053_ = new_n10051_;
  assign new_n10054_ = new_n4459_;
  assign new_n10055_ = new_n10054_;
  assign new_n10056_ = new_n10055_;
  assign new_n10057_ = new_n10055_;
  assign new_n10058_ = new_n10054_;
  assign new_n10059_ = new_n4458_;
  assign new_n10060_ = new_n10059_;
  assign new_n10061_ = new_n10060_;
  assign new_n10062_ = new_n10060_;
  assign new_n10063_ = new_n10059_;
  assign new_n10064_ = new_n10063_;
  assign new_n10065_ = new_n4521_;
  assign new_n10066_ = new_n4520_;
  assign new_n10067_ = new_n4463_;
  assign new_n10068_ = new_n10067_;
  assign new_n10069_ = new_n10068_;
  assign new_n10070_ = new_n10068_;
  assign new_n10071_ = new_n10067_;
  assign new_n10072_ = new_n4462_;
  assign new_n10073_ = new_n10072_;
  assign new_n10074_ = new_n10073_;
  assign new_n10075_ = new_n10073_;
  assign new_n10076_ = new_n10072_;
  assign new_n10077_ = new_n10076_;
  assign new_n10078_ = new_n4561_;
  assign new_n10079_ = new_n10078_;
  assign new_n10080_ = new_n10079_;
  assign new_n10081_ = new_n10079_;
  assign new_n10082_ = new_n10078_;
  assign new_n10083_ = new_n10082_;
  assign new_n10084_ = new_n10082_;
  assign new_n10085_ = new_n3951_;
  assign new_n10086_ = new_n4560_;
  assign new_n10087_ = new_n10086_;
  assign new_n10088_ = new_n10087_;
  assign new_n10089_ = new_n10088_;
  assign new_n10090_ = new_n10087_;
  assign new_n10091_ = new_n10086_;
  assign new_n10092_ = new_n10091_;
  assign new_n10093_ = new_n10091_;
  assign new_n10094_ = new_n3950_;
  assign new_n10095_ = new_n10094_;
  assign new_n10096_ = new_n10095_;
  assign new_n10097_ = new_n10094_;
  assign new_n10098_ = new_n4567_;
  assign new_n10099_ = new_n10098_;
  assign new_n10100_ = new_n10099_;
  assign new_n10101_ = new_n10099_;
  assign new_n10102_ = new_n10098_;
  assign new_n10103_ = new_n10102_;
  assign new_n10104_ = new_n10102_;
  assign new_n10105_ = new_n4566_;
  assign new_n10106_ = new_n10105_;
  assign new_n10107_ = new_n10106_;
  assign new_n10108_ = new_n10107_;
  assign new_n10109_ = new_n10106_;
  assign new_n10110_ = new_n10105_;
  assign new_n10111_ = new_n10110_;
  assign new_n10112_ = new_n10110_;
  assign new_n10113_ = new_n4517_;
  assign new_n10114_ = new_n4516_;
  assign new_n10115_ = new_n3927_;
  assign new_n10116_ = new_n3926_;
  assign new_n10117_ = new_n10116_;
  assign new_n10118_ = new_n10117_;
  assign new_n10119_ = new_n10116_;
  assign new_n10120_ = new_n6679_;
  assign new_n10121_ = new_n6658_;
  assign new_n10122_ = new_n6678_;
  assign new_n10123_ = new_n6659_;
  assign new_n10124_ = new_n4529_;
  assign new_n10125_ = new_n4528_;
  assign new_n10126_ = new_n3985_;
  assign new_n10127_ = new_n3984_;
  assign new_n10128_ = new_n10127_;
  assign new_n10129_ = new_n10128_;
  assign new_n10130_ = new_n10127_;
  assign new_n10131_ = new_n6704_;
  assign new_n10132_ = new_n6189_;
  assign new_n10133_ = new_n6705_;
  assign new_n10134_ = new_n6190_;
  assign new_n10135_ = new_n10134_;
  assign new_n10136_ = new_n4523_;
  assign new_n10137_ = new_n4522_;
  assign new_n10138_ = new_n3953_;
  assign new_n10139_ = new_n3952_;
  assign new_n10140_ = new_n10139_;
  assign new_n10141_ = new_n10140_;
  assign new_n10142_ = new_n10139_;
  assign new_n10143_ = new_n4519_;
  assign new_n10144_ = new_n4518_;
  assign new_n10145_ = new_n3931_;
  assign new_n10146_ = new_n3930_;
  assign new_n10147_ = new_n10146_;
  assign new_n10148_ = new_n10147_;
  assign new_n10149_ = new_n10146_;
  assign new_n10150_ = new_n6754_;
  assign new_n10151_ = new_n6733_;
  assign new_n10152_ = new_n6753_;
  assign new_n10153_ = new_n6734_;
  assign new_n10154_ = new_n4015_;
  assign new_n10155_ = new_n4014_;
  assign new_n10156_ = new_n10155_;
  assign new_n10157_ = new_n10156_;
  assign new_n10158_ = new_n10155_;
  assign new_n10159_ = new_n4243_;
  assign new_n10160_ = new_n4242_;
  assign new_n10161_ = new_n10160_;
  assign new_n10162_ = new_n10161_;
  assign new_n10163_ = new_n10160_;
  assign new_n10164_ = new_n6771_;
  assign new_n10165_ = new_n6765_;
  assign new_n10166_ = new_n6772_;
  assign new_n10167_ = new_n6766_;
  assign new_n10168_ = new_n4511_;
  assign new_n10169_ = new_n4510_;
  assign new_n10170_ = new_n4509_;
  assign new_n10171_ = new_n4508_;
  assign new_n10172_ = new_n6841_;
  assign new_n10173_ = new_n6820_;
  assign new_n10174_ = new_n6840_;
  assign new_n10175_ = new_n6821_;
  assign new_n10176_ = new_n6871_;
  assign new_n10177_ = new_n6858_;
  assign new_n10178_ = new_n6870_;
  assign new_n10179_ = new_n6859_;
  assign new_n10180_ = new_n6847_;
  assign new_n10181_ = new_n6800_;
  assign new_n10182_ = new_n6876_;
  assign new_n10183_ = new_n6801_;
  assign new_n10184_ = new_n6877_;
  assign new_n10185_ = new_n6846_;
  assign new_n10186_ = new_n4515_;
  assign new_n10187_ = new_n4514_;
  assign new_n10188_ = new_n4513_;
  assign new_n10189_ = new_n4512_;
  assign new_n10190_ = new_n6928_;
  assign new_n10191_ = new_n6907_;
  assign new_n10192_ = new_n6927_;
  assign new_n10193_ = new_n6908_;
  assign new_n10194_ = new_n6952_;
  assign new_n10195_ = new_n6939_;
  assign new_n10196_ = new_n6951_;
  assign new_n10197_ = new_n6940_;
  assign new_n10198_ = new_n6933_;
  assign new_n10199_ = new_n6272_;
  assign new_n10200_ = new_n6958_;
  assign new_n10201_ = new_n6271_;
  assign new_n10202_ = new_n10201_;
  assign new_n10203_ = new_n6957_;
  assign new_n10204_ = new_n6934_;
  assign new_n10205_ = new_n6553_;
  assign new_n10206_ = new_n10205_;
  assign new_n10207_ = new_n3558_;
  assign new_n10208_ = new_n10207_;
  assign new_n10209_ = new_n6547_;
  assign new_n10210_ = new_n10209_;
  assign new_n10211_ = new_n3586_;
  assign new_n10212_ = new_n10211_;
  assign new_n10213_ = new_n4540_;
  assign new_n10214_ = new_n6980_;
  assign new_n10215_ = new_n6979_;
  assign new_n10216_ = new_n6981_;
  assign new_n10217_ = new_n6978_;
  assign new_n10218_ = new_n6986_;
  assign new_n10219_ = new_n4157_;
  assign new_n10220_ = new_n10219_;
  assign new_n10221_ = new_n10219_;
  assign new_n10222_ = new_n6987_;
  assign new_n10223_ = new_n4156_;
  assign new_n10224_ = new_n10223_;
  assign new_n10225_ = new_n10224_;
  assign new_n10226_ = new_n10223_;
  assign new_n10227_ = new_n4140_;
  assign new_n10228_ = new_n10227_;
  assign new_n10229_ = new_n4141_;
  assign new_n10230_ = new_n4538_;
  assign new_n10231_ = new_n7005_;
  assign new_n10232_ = new_n7004_;
  assign new_n10233_ = new_n7006_;
  assign new_n10234_ = new_n7003_;
  assign new_n10235_ = new_n7011_;
  assign new_n10236_ = new_n4246_;
  assign new_n10237_ = new_n10236_;
  assign new_n10238_ = new_n10237_;
  assign new_n10239_ = new_n10236_;
  assign new_n10240_ = new_n7012_;
  assign new_n10241_ = new_n4247_;
  assign new_n10242_ = new_n10241_;
  assign new_n10243_ = new_n10241_;
  assign new_n10244_ = new_n4144_;
  assign new_n10245_ = new_n10244_;
  assign new_n10246_ = new_n4145_;
  assign new_n10247_ = new_n6280_;
  assign new_n10248_ = new_n10247_;
  assign new_n10249_ = new_n10247_;
  assign new_n10250_ = new_n4542_;
  assign new_n10251_ = new_n6279_;
  assign new_n10252_ = new_n10251_;
  assign new_n10253_ = new_n4488_;
  assign new_n10254_ = new_n10253_;
  assign new_n10255_ = new_n10254_;
  assign new_n10256_ = new_n10254_;
  assign new_n10257_ = new_n10253_;
  assign new_n10258_ = new_n10257_;
  assign new_n10259_ = new_n4454_;
  assign new_n10260_ = new_n10259_;
  assign new_n10261_ = new_n10259_;
  assign new_n10262_ = new_n4489_;
  assign new_n10263_ = new_n4455_;
  assign new_n10264_ = new_n10263_;
  assign new_n10265_ = new_n4612_;
  assign new_n10266_ = new_n10265_;
  assign new_n10267_ = new_n10265_;
  assign new_n10268_ = new_n4613_;
  assign new_n10269_ = new_n10268_;
  assign new_n10270_ = new_n6281_;
  assign new_n10271_ = new_n7034_;
  assign new_n10272_ = new_n10271_;
  assign new_n10273_ = new_n7035_;
  assign new_n10274_ = new_n10273_;
  assign new_n10275_ = new_n4659_;
  assign new_n10276_ = new_n10275_;
  assign new_n10277_ = new_n4658_;
  assign new_n10278_ = new_n10277_;
  assign new_n10279_ = new_n4240_;
  assign new_n10280_ = new_n4234_;
  assign new_n10281_ = new_n7041_;
  assign new_n10282_ = new_n7039_;
  assign new_n10283_ = new_n7040_;
  assign new_n10284_ = new_n7038_;
  assign new_n10285_ = new_n7046_;
  assign new_n10286_ = new_n7037_;
  assign new_n10287_ = new_n7047_;
  assign new_n10288_ = new_n7036_;
  assign new_n10289_ = new_n7061_;
  assign new_n10290_ = new_n7062_;
  assign new_n10291_ = new_n6273_;
  assign new_n10292_ = new_n10291_;
  assign new_n10293_ = new_n10291_;
  assign new_n10294_ = new_n4544_;
  assign new_n10295_ = new_n6274_;
  assign new_n10296_ = new_n10295_;
  assign new_n10297_ = new_n10296_;
  assign new_n10298_ = new_n10296_;
  assign new_n10299_ = new_n10295_;
  assign new_n10300_ = new_n10299_;
  assign new_n10301_ = new_n4490_;
  assign new_n10302_ = new_n10301_;
  assign new_n10303_ = new_n10302_;
  assign new_n10304_ = new_n10302_;
  assign new_n10305_ = new_n10301_;
  assign new_n10306_ = new_n10305_;
  assign new_n10307_ = new_n4456_;
  assign new_n10308_ = new_n10307_;
  assign new_n10309_ = new_n10307_;
  assign new_n10310_ = new_n4491_;
  assign new_n10311_ = new_n4457_;
  assign new_n10312_ = new_n10311_;
  assign new_n10313_ = new_n4614_;
  assign new_n10314_ = new_n10313_;
  assign new_n10315_ = new_n10313_;
  assign new_n10316_ = new_n4615_;
  assign new_n10317_ = new_n10316_;
  assign new_n10318_ = new_n7084_;
  assign new_n10319_ = new_n10318_;
  assign new_n10320_ = new_n7085_;
  assign new_n10321_ = new_n10320_;
  assign new_n10322_ = new_n4661_;
  assign new_n10323_ = new_n10322_;
  assign new_n10324_ = new_n4660_;
  assign new_n10325_ = new_n10324_;
  assign new_n10326_ = new_n4238_;
  assign new_n10327_ = new_n4236_;
  assign new_n10328_ = new_n7091_;
  assign new_n10329_ = new_n7089_;
  assign new_n10330_ = new_n7090_;
  assign new_n10331_ = new_n7088_;
  assign new_n10332_ = new_n7096_;
  assign new_n10333_ = new_n7087_;
  assign new_n10334_ = new_n7097_;
  assign new_n10335_ = new_n7086_;
  assign new_n10336_ = new_n7111_;
  assign new_n10337_ = new_n7112_;
  assign new_n10338_ = new_n3388_;
  assign new_n10339_ = new_n6359_;
  assign new_n10340_ = new_n10339_;
  assign new_n10341_ = new_n3596_;
  assign new_n10342_ = new_n10341_;
  assign new_n10343_ = new_n6360_;
  assign new_n10344_ = new_n10343_;
  assign new_n10345_ = new_n3597_;
  assign new_n10346_ = new_n10345_;
  assign new_n10347_ = new_n3550_;
  assign new_n10348_ = new_n10347_;
  assign new_n10349_ = new_n6366_;
  assign new_n10350_ = new_n10349_;
  assign new_n10351_ = new_n3578_;
  assign new_n10352_ = new_n10351_;
  assign new_n10353_ = new_n6378_;
  assign new_n10354_ = new_n10353_;
  assign new_n10355_ = new_n3582_;
  assign new_n10356_ = new_n10355_;
  assign new_n10357_ = new_n6372_;
  assign new_n10358_ = new_n10357_;
  assign new_n10359_ = new_n4160_;
  assign new_n10360_ = new_n10359_;
  assign new_n10361_ = new_n3431_;
  assign new_n10362_ = new_n10361_;
  assign new_n10363_ = new_n3435_;
  assign new_n10364_ = new_n10363_;
  assign new_n10365_ = new_n4128_;
  assign new_n10366_ = new_n10365_;
  assign new_n10367_ = new_n10365_;
  assign new_n10368_ = new_n6535_;
  assign new_n10369_ = new_n10368_;
  assign new_n10370_ = new_n3571_;
  assign new_n10371_ = new_n4662_;
  assign new_n10372_ = new_n4655_;
  assign new_n10373_ = new_n4663_;
  assign new_n10374_ = new_n4654_;
  assign new_n10375_ = new_n7161_;
  assign new_n10376_ = new_n7162_;
  assign new_n10377_ = new_n7171_;
  assign new_n10378_ = new_n6538_;
  assign new_n10379_ = new_n10378_;
  assign new_n10380_ = new_n10379_;
  assign new_n10381_ = new_n10378_;
  assign new_n10382_ = new_n4665_;
  assign new_n10383_ = new_n4657_;
  assign new_n10384_ = new_n4664_;
  assign new_n10385_ = new_n4656_;
  assign new_n10386_ = new_n7177_;
  assign new_n10387_ = new_n7178_;
  assign new_n10388_ = new_n7187_;
  assign new_n10389_ = new_n6541_;
  assign new_n10390_ = new_n10389_;
  assign new_n10391_ = new_n10390_;
  assign new_n10392_ = new_n10389_;
  assign new_n10393_ = new_n3466_;
  assign new_n10394_ = new_n3472_;
  assign new_n10395_ = new_n6328_;
  assign new_n10396_ = new_n10395_;
  assign new_n10397_ = new_n10395_;
  assign new_n10398_ = new_n6305_;
  assign new_n10399_ = new_n10398_;
  assign new_n10400_ = new_n6327_;
  assign new_n10401_ = new_n10400_;
  assign new_n10402_ = new_n6306_;
  assign new_n10403_ = new_n7202_;
  assign new_n10404_ = new_n7133_;
  assign new_n10405_ = new_n10404_;
  assign new_n10406_ = new_n10405_;
  assign new_n10407_ = new_n10404_;
  assign new_n10408_ = new_n6340_;
  assign new_n10409_ = new_n10408_;
  assign new_n10410_ = new_n6307_;
  assign new_n10411_ = new_n10410_;
  assign new_n10412_ = new_n6339_;
  assign new_n10413_ = new_n10412_;
  assign new_n10414_ = new_n6308_;
  assign new_n10415_ = new_n7206_;
  assign new_n10416_ = new_n7129_;
  assign new_n10417_ = new_n10416_;
  assign new_n10418_ = new_n10416_;
  assign new_n10419_ = new_n6334_;
  assign new_n10420_ = new_n10419_;
  assign new_n10421_ = new_n10420_;
  assign new_n10422_ = new_n10420_;
  assign new_n10423_ = new_n10419_;
  assign new_n10424_ = new_n6333_;
  assign new_n10425_ = new_n10424_;
  assign new_n10426_ = new_n6321_;
  assign new_n10427_ = new_n10426_;
  assign new_n10428_ = new_n10427_;
  assign new_n10429_ = new_n10426_;
  assign new_n10430_ = new_n6322_;
  assign new_n10431_ = new_n10430_;
  assign new_n10432_ = new_n10430_;
  assign new_n10433_ = new_n7210_;
  assign new_n10434_ = new_n3476_;
  assign new_n10435_ = new_n6356_;
  assign new_n10436_ = new_n10435_;
  assign new_n10437_ = new_n7214_;
  assign new_n10438_ = new_n6346_;
  assign new_n10439_ = new_n10438_;
  assign new_n10440_ = new_n6345_;
  assign new_n10441_ = new_n10440_;
  assign new_n10442_ = new_n10440_;
  assign new_n10443_ = new_n6299_;
  assign new_n10444_ = new_n10443_;
  assign new_n10445_ = new_n10443_;
  assign new_n10446_ = new_n6300_;
  assign new_n10447_ = new_n10446_;
  assign new_n10448_ = new_n10447_;
  assign new_n10449_ = new_n10447_;
  assign new_n10450_ = new_n10446_;
  assign new_n10451_ = new_n10450_;
  assign new_n10452_ = new_n10450_;
  assign new_n10453_ = new_n7221_;
  assign new_n10454_ = new_n7223_;
  assign new_n10455_ = new_n6347_;
  assign new_n10456_ = new_n10455_;
  assign new_n10457_ = new_n6350_;
  assign new_n10458_ = new_n6349_;
  assign new_n10459_ = new_n7231_;
  assign new_n10460_ = new_n10459_;
  assign new_n10461_ = new_n7234_;
  assign new_n10462_ = new_n7237_;
  assign new_n10463_ = new_n7238_;
  assign new_n10464_ = new_n7233_;
  assign new_n10465_ = new_n7243_;
  assign new_n10466_ = new_n7250_;
  assign new_n10467_ = new_n10466_;
  assign new_n10468_ = new_n7251_;
  assign new_n10469_ = new_n10468_;
  assign new_n10470_ = new_n7258_;
  assign new_n10471_ = new_n7245_;
  assign new_n10472_ = new_n7197_;
  assign new_n10473_ = new_n7136_;
  assign new_n10474_ = new_n10473_;
  assign new_n10475_ = new_n7200_;
  assign new_n10476_ = new_n7139_;
  assign new_n10477_ = new_n10476_;
  assign new_n10478_ = new_n7226_;
  assign new_n10479_ = new_n7153_;
  assign new_n10480_ = new_n7204_;
  assign new_n10481_ = new_n7212_;
  assign new_n10482_ = new_n7227_;
  assign new_n10483_ = new_n7152_;
  assign new_n10484_ = new_n7207_;
  assign new_n10485_ = new_n7222_;
  assign new_n10486_ = new_n6970_;
  assign new_n10487_ = new_n7154_;
  assign new_n10488_ = new_n6971_;
  assign new_n10489_ = new_n7155_;
  assign new_n10490_ = new_n7232_;
  assign new_n10491_ = new_n2578_;
  assign new_n10492_ = new_n2572_;
  assign new_n10493_ = new_n10492_;
  assign new_n10494_ = new_n10493_;
  assign new_n10495_ = new_n10492_;
  assign new_n10496_ = new_n2580_;
  assign new_n10497_ = new_n2573_;
  assign new_n10498_ = new_n2582_;
  assign new_n10499_ = new_n2584_;
  assign new_n10500_ = new_n2574_;
  assign new_n10501_ = new_n10500_;
  assign new_n10502_ = new_n10501_;
  assign new_n10503_ = new_n10501_;
  assign new_n10504_ = new_n10500_;
  assign new_n10505_ = new_n2536_;
  assign new_n10506_ = new_n2575_;
  assign new_n10507_ = new_n10506_;
  assign new_n10508_ = new_n2540_;
  assign new_n10509_ = new_n2544_;
  assign new_n10510_ = new_n3611_;
  assign new_n10511_ = new_n10510_;
  assign new_n10512_ = new_n3618_;
  assign new_n10513_ = new_n2691_;
  assign new_n10514_ = new_n10513_;
  assign new_n10515_ = new_n10513_;
  assign new_n10516_ = new_n3475_;
  assign new_n10517_ = new_n4726_;
  assign new_n10518_ = new_n4038_;
  assign new_n10519_ = new_n4248_;
  assign new_n10520_ = new_n10519_;
  assign new_n10521_ = new_n4044_;
  assign new_n10522_ = new_n10521_;
  assign new_n10523_ = new_n10521_;
  assign new_n10524_ = new_n4046_;
  assign new_n10525_ = new_n10524_;
  assign new_n10526_ = new_n10524_;
  assign new_n10527_ = new_n4048_;
  assign new_n10528_ = new_n10527_;
  assign new_n10529_ = new_n10527_;
  assign new_n10530_ = new_n4052_;
  assign new_n10531_ = new_n10530_;
  assign new_n10532_ = new_n10530_;
  assign new_n10533_ = new_n4126_;
  assign new_n10534_ = new_n4130_;
  assign new_n10535_ = new_n4152_;
  assign new_n10536_ = new_n4154_;
  assign new_n10537_ = new_n4250_;
  assign new_n10538_ = new_n6422_;
  assign new_n10539_ = new_n6451_;
  assign new_n10540_ = new_n6494_;
  assign new_n10541_ = new_n6523_;
  assign new_n10542_ = new_n6529_;
  assign new_n10543_ = new_n3430_;
  assign new_n10544_ = new_n3434_;
  assign new_n10545_ = new_n6996_;
  assign new_n10546_ = new_n7021_;
  assign new_n10547_ = new_n7056_;
  assign new_n10548_ = new_n7071_;
  assign new_n10549_ = new_n7106_;
  assign new_n10550_ = new_n7121_;
  assign new_n10551_ = new_n3574_;
  assign new_n10552_ = new_n10551_;
  assign new_n10553_ = new_n7124_;
  assign new_n10554_ = new_n10553_;
  assign new_n10555_ = new_n3418_;
  assign new_n10556_ = new_n3438_;
  assign new_n10557_ = new_n7294_;
  assign new_n10558_ = new_n7297_;
  assign new_n10559_ = new_n7300_;
  assign new_n10560_ = new_n7303_;
  assign new_n10561_ = new_n2602_;
  assign new_n10562_ = new_n2604_;
  assign new_n10563_ = new_n2624_;
  assign new_n10564_ = new_n2626_;
  always @ (posedge clock) begin
    n2610_lo <= n2610_li;
    n2613_lo <= n2613_li;
    n2616_lo <= n2616_li;
    n2619_lo <= n2619_li;
    n2622_lo <= n2622_li;
    n2625_lo <= n2625_li;
    n2628_lo <= n2628_li;
    n2631_lo <= n2631_li;
    n2634_lo <= n2634_li;
    n2637_lo <= n2637_li;
    n2640_lo <= n2640_li;
    n2643_lo <= n2643_li;
    n2646_lo <= n2646_li;
    n2649_lo <= n2649_li;
    n2652_lo <= n2652_li;
    n2655_lo <= n2655_li;
    n2658_lo <= n2658_li;
    n2661_lo <= n2661_li;
    n2664_lo <= n2664_li;
    n2667_lo <= n2667_li;
    n2670_lo <= n2670_li;
    n2673_lo <= n2673_li;
    n2676_lo <= n2676_li;
    n2679_lo <= n2679_li;
    n2682_lo <= n2682_li;
    n2685_lo <= n2685_li;
    n2688_lo <= n2688_li;
    n2691_lo <= n2691_li;
    n2694_lo <= n2694_li;
    n2697_lo <= n2697_li;
    n2700_lo <= n2700_li;
    n2703_lo <= n2703_li;
    n2706_lo <= n2706_li;
    n2709_lo <= n2709_li;
    n2712_lo <= n2712_li;
    n2715_lo <= n2715_li;
    n2718_lo <= n2718_li;
    n2721_lo <= n2721_li;
    n2724_lo <= n2724_li;
    n2727_lo <= n2727_li;
    n2730_lo <= n2730_li;
    n2733_lo <= n2733_li;
    n2736_lo <= n2736_li;
    n2739_lo <= n2739_li;
    n2742_lo <= n2742_li;
    n2745_lo <= n2745_li;
    n2748_lo <= n2748_li;
    n2751_lo <= n2751_li;
    n2754_lo <= n2754_li;
    n2757_lo <= n2757_li;
    n2760_lo <= n2760_li;
    n2763_lo <= n2763_li;
    n2766_lo <= n2766_li;
    n2769_lo <= n2769_li;
    n2772_lo <= n2772_li;
    n2775_lo <= n2775_li;
    n2778_lo <= n2778_li;
    n2781_lo <= n2781_li;
    n2784_lo <= n2784_li;
    n2787_lo <= n2787_li;
    n2790_lo <= n2790_li;
    n2793_lo <= n2793_li;
    n2796_lo <= n2796_li;
    n2799_lo <= n2799_li;
    n2802_lo <= n2802_li;
    n2805_lo <= n2805_li;
    n2808_lo <= n2808_li;
    n2811_lo <= n2811_li;
    n2814_lo <= n2814_li;
    n2817_lo <= n2817_li;
    n2820_lo <= n2820_li;
    n2823_lo <= n2823_li;
    n2826_lo <= n2826_li;
    n2829_lo <= n2829_li;
    n2832_lo <= n2832_li;
    n2835_lo <= n2835_li;
    n2838_lo <= n2838_li;
    n2841_lo <= n2841_li;
    n2844_lo <= n2844_li;
    n2847_lo <= n2847_li;
    n2850_lo <= n2850_li;
    n2853_lo <= n2853_li;
    n2856_lo <= n2856_li;
    n2859_lo <= n2859_li;
    n2862_lo <= n2862_li;
    n2865_lo <= n2865_li;
    n2868_lo <= n2868_li;
    n2871_lo <= n2871_li;
    n2874_lo <= n2874_li;
    n2877_lo <= n2877_li;
    n2880_lo <= n2880_li;
    n2883_lo <= n2883_li;
    n2886_lo <= n2886_li;
    n2889_lo <= n2889_li;
    n2892_lo <= n2892_li;
    n2895_lo <= n2895_li;
    n2898_lo <= n2898_li;
    n2901_lo <= n2901_li;
    n2904_lo <= n2904_li;
    n2907_lo <= n2907_li;
    n2910_lo <= n2910_li;
    n2913_lo <= n2913_li;
    n2916_lo <= n2916_li;
    n2919_lo <= n2919_li;
    n2922_lo <= n2922_li;
    n2925_lo <= n2925_li;
    n2928_lo <= n2928_li;
    n2931_lo <= n2931_li;
    n2934_lo <= n2934_li;
    n2937_lo <= n2937_li;
    n2940_lo <= n2940_li;
    n2943_lo <= n2943_li;
    n2946_lo <= n2946_li;
    n2949_lo <= n2949_li;
    n2952_lo <= n2952_li;
    n2955_lo <= n2955_li;
    n2958_lo <= n2958_li;
    n2961_lo <= n2961_li;
    n2964_lo <= n2964_li;
    n2967_lo <= n2967_li;
    n2970_lo <= n2970_li;
    n2973_lo <= n2973_li;
    n2976_lo <= n2976_li;
    n2979_lo <= n2979_li;
    n2982_lo <= n2982_li;
    n2985_lo <= n2985_li;
    n2988_lo <= n2988_li;
    n2991_lo <= n2991_li;
    n2994_lo <= n2994_li;
    n2997_lo <= n2997_li;
    n3000_lo <= n3000_li;
    n3003_lo <= n3003_li;
    n3006_lo <= n3006_li;
    n3009_lo <= n3009_li;
    n3012_lo <= n3012_li;
    n3015_lo <= n3015_li;
    n3018_lo <= n3018_li;
    n3021_lo <= n3021_li;
    n3024_lo <= n3024_li;
    n3027_lo <= n3027_li;
    n3030_lo <= n3030_li;
    n3033_lo <= n3033_li;
    n3036_lo <= n3036_li;
    n3039_lo <= n3039_li;
    n3042_lo <= n3042_li;
    n3045_lo <= n3045_li;
    n3048_lo <= n3048_li;
    n3051_lo <= n3051_li;
    n3054_lo <= n3054_li;
    n3057_lo <= n3057_li;
    n3060_lo <= n3060_li;
    n3063_lo <= n3063_li;
    n3066_lo <= n3066_li;
    n3069_lo <= n3069_li;
    n3072_lo <= n3072_li;
    n3075_lo <= n3075_li;
    n3078_lo <= n3078_li;
    n3081_lo <= n3081_li;
    n3084_lo <= n3084_li;
    n3087_lo <= n3087_li;
    n3090_lo <= n3090_li;
    n3093_lo <= n3093_li;
    n3096_lo <= n3096_li;
    n3099_lo <= n3099_li;
    n3102_lo <= n3102_li;
    n3105_lo <= n3105_li;
    n3108_lo <= n3108_li;
    n3111_lo <= n3111_li;
    n3114_lo <= n3114_li;
    n3117_lo <= n3117_li;
    n3120_lo <= n3120_li;
    n3123_lo <= n3123_li;
    n3126_lo <= n3126_li;
    n3129_lo <= n3129_li;
    n3132_lo <= n3132_li;
    n3135_lo <= n3135_li;
    n3138_lo <= n3138_li;
    n3141_lo <= n3141_li;
    n3144_lo <= n3144_li;
    n3147_lo <= n3147_li;
    n3150_lo <= n3150_li;
    n3153_lo <= n3153_li;
    n3156_lo <= n3156_li;
    n3159_lo <= n3159_li;
    n3162_lo <= n3162_li;
    n3165_lo <= n3165_li;
    n3168_lo <= n3168_li;
    n3171_lo <= n3171_li;
    n3174_lo <= n3174_li;
    n3177_lo <= n3177_li;
    n3180_lo <= n3180_li;
    n3183_lo <= n3183_li;
    n3186_lo <= n3186_li;
    n3189_lo <= n3189_li;
    n3192_lo <= n3192_li;
    n3195_lo <= n3195_li;
    n3198_lo <= n3198_li;
    n3201_lo <= n3201_li;
    n3204_lo <= n3204_li;
    n3207_lo <= n3207_li;
    n3210_lo <= n3210_li;
    n3213_lo <= n3213_li;
    n3216_lo <= n3216_li;
    n3219_lo <= n3219_li;
    n3222_lo <= n3222_li;
    n3225_lo <= n3225_li;
    n3228_lo <= n3228_li;
    n3231_lo <= n3231_li;
    n3234_lo <= n3234_li;
    n3237_lo <= n3237_li;
    n3240_lo <= n3240_li;
    n3243_lo <= n3243_li;
    n3246_lo <= n3246_li;
    n3249_lo <= n3249_li;
    n3252_lo <= n3252_li;
    n3255_lo <= n3255_li;
    n3258_lo <= n3258_li;
    n3261_lo <= n3261_li;
    n3264_lo <= n3264_li;
    n3267_lo <= n3267_li;
    n3270_lo <= n3270_li;
    n3273_lo <= n3273_li;
    n3276_lo <= n3276_li;
    n3279_lo <= n3279_li;
    n3282_lo <= n3282_li;
    n3285_lo <= n3285_li;
    n3288_lo <= n3288_li;
    n3291_lo <= n3291_li;
    n3294_lo <= n3294_li;
    n3297_lo <= n3297_li;
    n3300_lo <= n3300_li;
    n3303_lo <= n3303_li;
    n3306_lo <= n3306_li;
    n3309_lo <= n3309_li;
    n3312_lo <= n3312_li;
    n3315_lo <= n3315_li;
    n3318_lo <= n3318_li;
    n3321_lo <= n3321_li;
    n3324_lo <= n3324_li;
    n3327_lo <= n3327_li;
    n3330_lo <= n3330_li;
    n3333_lo <= n3333_li;
    n3336_lo <= n3336_li;
    n3339_lo <= n3339_li;
    n3342_lo <= n3342_li;
    n3345_lo <= n3345_li;
    n3348_lo <= n3348_li;
    n3351_lo <= n3351_li;
    n3354_lo <= n3354_li;
    n3357_lo <= n3357_li;
    n3360_lo <= n3360_li;
    n3363_lo <= n3363_li;
    n3366_lo <= n3366_li;
    n3369_lo <= n3369_li;
    n3372_lo <= n3372_li;
    n3375_lo <= n3375_li;
    n3378_lo <= n3378_li;
    n3381_lo <= n3381_li;
    n3384_lo <= n3384_li;
    n3387_lo <= n3387_li;
    n3390_lo <= n3390_li;
    n3393_lo <= n3393_li;
    n3396_lo <= n3396_li;
    n3399_lo <= n3399_li;
    n3402_lo <= n3402_li;
    n3405_lo <= n3405_li;
    n3408_lo <= n3408_li;
    n3411_lo <= n3411_li;
    n3414_lo <= n3414_li;
    n3417_lo <= n3417_li;
    n3420_lo <= n3420_li;
    n3423_lo <= n3423_li;
    n3426_lo <= n3426_li;
    n3429_lo <= n3429_li;
    n3432_lo <= n3432_li;
    n3435_lo <= n3435_li;
    n3438_lo <= n3438_li;
    n3441_lo <= n3441_li;
    n3444_lo <= n3444_li;
    n3447_lo <= n3447_li;
    n3450_lo <= n3450_li;
    n3453_lo <= n3453_li;
    n3456_lo <= n3456_li;
    n3459_lo <= n3459_li;
    n3462_lo <= n3462_li;
    n3465_lo <= n3465_li;
    n3468_lo <= n3468_li;
    n3471_lo <= n3471_li;
    n3474_lo <= n3474_li;
    n3477_lo <= n3477_li;
    n3480_lo <= n3480_li;
    n3483_lo <= n3483_li;
    n3486_lo <= n3486_li;
    n3489_lo <= n3489_li;
    n3492_lo <= n3492_li;
    n3495_lo <= n3495_li;
    n3498_lo <= n3498_li;
    n3501_lo <= n3501_li;
    n3504_lo <= n3504_li;
    n3507_lo <= n3507_li;
    n3510_lo <= n3510_li;
    n3513_lo <= n3513_li;
    n3516_lo <= n3516_li;
    n3519_lo <= n3519_li;
    n3522_lo <= n3522_li;
    n3525_lo <= n3525_li;
    n3528_lo <= n3528_li;
    n3531_lo <= n3531_li;
    n3534_lo <= n3534_li;
    n3537_lo <= n3537_li;
    n3540_lo <= n3540_li;
    n3543_lo <= n3543_li;
    n3546_lo <= n3546_li;
    n3549_lo <= n3549_li;
    n3552_lo <= n3552_li;
    n3555_lo <= n3555_li;
    n3558_lo <= n3558_li;
    n3561_lo <= n3561_li;
    n3564_lo <= n3564_li;
    n3567_lo <= n3567_li;
    n3570_lo <= n3570_li;
    n3573_lo <= n3573_li;
    n3576_lo <= n3576_li;
    n3579_lo <= n3579_li;
    n3582_lo <= n3582_li;
    n3585_lo <= n3585_li;
    n3588_lo <= n3588_li;
    n3591_lo <= n3591_li;
    n3594_lo <= n3594_li;
    n3597_lo <= n3597_li;
    n3600_lo <= n3600_li;
    n3603_lo <= n3603_li;
    n3606_lo <= n3606_li;
    n3609_lo <= n3609_li;
    n3612_lo <= n3612_li;
    n3615_lo <= n3615_li;
    n3618_lo <= n3618_li;
    n3621_lo <= n3621_li;
    n3624_lo <= n3624_li;
    n3627_lo <= n3627_li;
    n3630_lo <= n3630_li;
    n3633_lo <= n3633_li;
    n3636_lo <= n3636_li;
    n3639_lo <= n3639_li;
    n3642_lo <= n3642_li;
    n3645_lo <= n3645_li;
    n3648_lo <= n3648_li;
    n3651_lo <= n3651_li;
    n3654_lo <= n3654_li;
    n3657_lo <= n3657_li;
    n3666_lo <= n3666_li;
    n3669_lo <= n3669_li;
    n3678_lo <= n3678_li;
    n3687_lo <= n3687_li;
    n3690_lo <= n3690_li;
    n3702_lo <= n3702_li;
    n3711_lo <= n3711_li;
    n3714_lo <= n3714_li;
    n3726_lo <= n3726_li;
    n3735_lo <= n3735_li;
    n3738_lo <= n3738_li;
    n3750_lo <= n3750_li;
    n3753_lo <= n3753_li;
    n3759_lo <= n3759_li;
    n3762_lo <= n3762_li;
    n3765_lo <= n3765_li;
    n3774_lo <= n3774_li;
    n3777_lo <= n3777_li;
    n3786_lo <= n3786_li;
    n3789_lo <= n3789_li;
    n3792_lo <= n3792_li;
    n3795_lo <= n3795_li;
    n3798_lo <= n3798_li;
    n3801_lo <= n3801_li;
    n3810_lo <= n3810_li;
    n3813_lo <= n3813_li;
    n3822_lo <= n3822_li;
    n3825_lo <= n3825_li;
    n3834_lo <= n3834_li;
    n3843_lo <= n3843_li;
    n3846_lo <= n3846_li;
    n3867_lo <= n3867_li;
    n3891_lo <= n3891_li;
    n3915_lo <= n3915_li;
    n3930_lo <= n3930_li;
    n3933_lo <= n3933_li;
    n3936_lo <= n3936_li;
    n3942_lo <= n3942_li;
    n3945_lo <= n3945_li;
    n3948_lo <= n3948_li;
    n3954_lo <= n3954_li;
    n3957_lo <= n3957_li;
    n3963_lo <= n3963_li;
    n3966_lo <= n3966_li;
    n3969_lo <= n3969_li;
    n3975_lo <= n3975_li;
    n3978_lo <= n3978_li;
    n3987_lo <= n3987_li;
    n3990_lo <= n3990_li;
    n4002_lo <= n4002_li;
    n4011_lo <= n4011_li;
    n4014_lo <= n4014_li;
    n4026_lo <= n4026_li;
    n4035_lo <= n4035_li;
    n4038_lo <= n4038_li;
    n4050_lo <= n4050_li;
    n4053_lo <= n4053_li;
    n4059_lo <= n4059_li;
    n4062_lo <= n4062_li;
    n4065_lo <= n4065_li;
    n4098_lo <= n4098_li;
    n4107_lo <= n4107_li;
    n4119_lo <= n4119_li;
    n4131_lo <= n4131_li;
    n4143_lo <= n4143_li;
    n4155_lo <= n4155_li;
    n4167_lo <= n4167_li;
    n4179_lo <= n4179_li;
    n4182_lo <= n4182_li;
    n4185_lo <= n4185_li;
    n4188_lo <= n4188_li;
    n4194_lo <= n4194_li;
    n4197_lo <= n4197_li;
    n4200_lo <= n4200_li;
    n4206_lo <= n4206_li;
    n4209_lo <= n4209_li;
    n4212_lo <= n4212_li;
    n4215_lo <= n4215_li;
    n4227_lo <= n4227_li;
    n4230_lo <= n4230_li;
    n4233_lo <= n4233_li;
    n4236_lo <= n4236_li;
    n4239_lo <= n4239_li;
    n4242_lo <= n4242_li;
    n4251_lo <= n4251_li;
    n4263_lo <= n4263_li;
    n4275_lo <= n4275_li;
    n4278_lo <= n4278_li;
    n4287_lo <= n4287_li;
    n4290_lo <= n4290_li;
    n4293_lo <= n4293_li;
    n4299_lo <= n4299_li;
    n4302_lo <= n4302_li;
    n4305_lo <= n4305_li;
    n4311_lo <= n4311_li;
    n4314_lo <= n4314_li;
    n4323_lo <= n4323_li;
    n4326_lo <= n4326_li;
    n4335_lo <= n4335_li;
    n4338_lo <= n4338_li;
    n4347_lo <= n4347_li;
    n4350_lo <= n4350_li;
    n4359_lo <= n4359_li;
    n4362_lo <= n4362_li;
    n4365_lo <= n4365_li;
    n4371_lo <= n4371_li;
    n4374_lo <= n4374_li;
    n4383_lo <= n4383_li;
    n4395_lo <= n4395_li;
    n4407_lo <= n4407_li;
    n4410_lo <= n4410_li;
    n4413_lo <= n4413_li;
    n4416_lo <= n4416_li;
    n4419_lo <= n4419_li;
    n4422_lo <= n4422_li;
    n4425_lo <= n4425_li;
    n4428_lo <= n4428_li;
    n4431_lo <= n4431_li;
    n4434_lo <= n4434_li;
    n4437_lo <= n4437_li;
    n4440_lo <= n4440_li;
    n4443_lo <= n4443_li;
    n4446_lo <= n4446_li;
    n4449_lo <= n4449_li;
    n4452_lo <= n4452_li;
    n4455_lo <= n4455_li;
    n4458_lo <= n4458_li;
    n4461_lo <= n4461_li;
    n4464_lo <= n4464_li;
    n4467_lo <= n4467_li;
    n4470_lo <= n4470_li;
    n4473_lo <= n4473_li;
    n4476_lo <= n4476_li;
    n4479_lo <= n4479_li;
    n4482_lo <= n4482_li;
    n4485_lo <= n4485_li;
    n4488_lo <= n4488_li;
    n4494_lo <= n4494_li;
    n4497_lo <= n4497_li;
    n4500_lo <= n4500_li;
    n4503_lo <= n4503_li;
    n4506_lo <= n4506_li;
    n4509_lo <= n4509_li;
    n4512_lo <= n4512_li;
    n4515_lo <= n4515_li;
    n4518_lo <= n4518_li;
    n4521_lo <= n4521_li;
    n4524_lo <= n4524_li;
    n4527_lo <= n4527_li;
    n4530_lo <= n4530_li;
    n4533_lo <= n4533_li;
    n4536_lo <= n4536_li;
    n4539_lo <= n4539_li;
    n4542_lo <= n4542_li;
    n4545_lo <= n4545_li;
    n4548_lo <= n4548_li;
    n4554_lo <= n4554_li;
    n4557_lo <= n4557_li;
    n4560_lo <= n4560_li;
    n4563_lo <= n4563_li;
    n4566_lo <= n4566_li;
    n4569_lo <= n4569_li;
    n4572_lo <= n4572_li;
    n4575_lo <= n4575_li;
    n4578_lo <= n4578_li;
    n4581_lo <= n4581_li;
    n4584_lo <= n4584_li;
    n4587_lo <= n4587_li;
    n4590_lo <= n4590_li;
    n4593_lo <= n4593_li;
    n4596_lo <= n4596_li;
    n4599_lo <= n4599_li;
    n4602_lo <= n4602_li;
    n4605_lo <= n4605_li;
    n4608_lo <= n4608_li;
    n4611_lo <= n4611_li;
    n4614_lo <= n4614_li;
    n4617_lo <= n4617_li;
    n4620_lo <= n4620_li;
    n4623_lo <= n4623_li;
    n4626_lo <= n4626_li;
    n4629_lo <= n4629_li;
    n4632_lo <= n4632_li;
    n4635_lo <= n4635_li;
    n4638_lo <= n4638_li;
    n4641_lo <= n4641_li;
    n4644_lo <= n4644_li;
    n4647_lo <= n4647_li;
    n4650_lo <= n4650_li;
    n4653_lo <= n4653_li;
    n4656_lo <= n4656_li;
    n4659_lo <= n4659_li;
    n4662_lo <= n4662_li;
    n4665_lo <= n4665_li;
    n4668_lo <= n4668_li;
    n4671_lo <= n4671_li;
    n4674_lo <= n4674_li;
    n4677_lo <= n4677_li;
    n4680_lo <= n4680_li;
    n4683_lo <= n4683_li;
    n4686_lo <= n4686_li;
    n4689_lo <= n4689_li;
    n4692_lo <= n4692_li;
    n4695_lo <= n4695_li;
    n4698_lo <= n4698_li;
    n4701_lo <= n4701_li;
    n4704_lo <= n4704_li;
    n4707_lo <= n4707_li;
    n4710_lo <= n4710_li;
    n4713_lo <= n4713_li;
    n4716_lo <= n4716_li;
    n4719_lo <= n4719_li;
    n4722_lo <= n4722_li;
    n4725_lo <= n4725_li;
    n4728_lo <= n4728_li;
    n4731_lo <= n4731_li;
    n4734_lo <= n4734_li;
    n4737_lo <= n4737_li;
    n4740_lo <= n4740_li;
    n4743_lo <= n4743_li;
    n6382_o2 <= n6382_i2;
    n6383_o2 <= n6383_i2;
    n6419_o2 <= n6419_i2;
    n6420_o2 <= n6420_i2;
    n6435_o2 <= n6435_i2;
    n6436_o2 <= n6436_i2;
    n6448_o2 <= n6448_i2;
    n6449_o2 <= n6449_i2;
    n6613_o2 <= n6613_i2;
    n6614_o2 <= n6614_i2;
    n6641_o2 <= n6641_i2;
    n6658_o2 <= n6658_i2;
    n6757_o2 <= n6757_i2;
    n6756_o2 <= n6756_i2;
    n7116_o2 <= n7116_i2;
    n7156_o2 <= n7156_i2;
    n6549_o2 <= n6549_i2;
    n6550_o2 <= n6550_i2;
    n7357_o2 <= n7357_i2;
    n7358_o2 <= n7358_i2;
    n7359_o2 <= n7359_i2;
    n7360_o2 <= n7360_i2;
    n6621_o2 <= n6621_i2;
    n6623_o2 <= n6623_i2;
    n6625_o2 <= n6625_i2;
    n6626_o2 <= n6626_i2;
    n6627_o2 <= n6627_i2;
    n6628_o2 <= n6628_i2;
    n6629_o2 <= n6629_i2;
    n6630_o2 <= n6630_i2;
    n6669_o2 <= n6669_i2;
    n7449_o2 <= n7449_i2;
    n7450_o2 <= n7450_i2;
    n7451_o2 <= n7451_i2;
    n7452_o2 <= n7452_i2;
    n6682_o2 <= n6682_i2;
    n6683_o2 <= n6683_i2;
    n6684_o2 <= n6684_i2;
    n6685_o2 <= n6685_i2;
    n7463_o2 <= n7463_i2;
    n6686_o2 <= n6686_i2;
    n6687_o2 <= n6687_i2;
    n6688_o2 <= n6688_i2;
    n6689_o2 <= n6689_i2;
    n6772_o2 <= n6772_i2;
    n6773_o2 <= n6773_i2;
    n6774_o2 <= n6774_i2;
    n6775_o2 <= n6775_i2;
    G3467_o2 <= G3467_i2;
    G2810_o2 <= G2810_i2;
    n6833_o2 <= n6833_i2;
    n6945_o2 <= n6945_i2;
    n6947_o2 <= n6947_i2;
    n6949_o2 <= n6949_i2;
    n6951_o2 <= n6951_i2;
    n6888_o2 <= n6888_i2;
    n6889_o2 <= n6889_i2;
    n6936_o2 <= n6936_i2;
    n6954_o2 <= n6954_i2;
    n6955_o2 <= n6955_i2;
    n6956_o2 <= n6956_i2;
    n6957_o2 <= n6957_i2;
    n6958_o2 <= n6958_i2;
    n6982_o2 <= n6982_i2;
    n6984_o2 <= n6984_i2;
    n6974_o2 <= n6974_i2;
    n6975_o2 <= n6975_i2;
    n6999_o2 <= n6999_i2;
    n7015_o2 <= n7015_i2;
    n7016_o2 <= n7016_i2;
    n7017_o2 <= n7017_i2;
    n7018_o2 <= n7018_i2;
    n7005_o2 <= n7005_i2;
    n7019_o2 <= n7019_i2;
    n7022_o2 <= n7022_i2;
    n7023_o2 <= n7023_i2;
    n7132_o2 <= n7132_i2;
    n7133_o2 <= n7133_i2;
    n7135_o2 <= n7135_i2;
    n7136_o2 <= n7136_i2;
    n7175_o2 <= n7175_i2;
    n7155_o2 <= n7155_i2;
    G3060_o2 <= G3060_i2;
    n7383_o2 <= n7383_i2;
    G3802_o2 <= G3802_i2;
    G3859_o2 <= G3859_i2;
    n7355_o2 <= n7355_i2;
    n7356_o2 <= n7356_i2;
    G4054_o2 <= G4054_i2;
    G4068_o2 <= G4068_i2;
    n7384_o2 <= n7384_i2;
    n7387_o2 <= n7387_i2;
    n7388_o2 <= n7388_i2;
    n7389_o2 <= n7389_i2;
    n7386_o2 <= n7386_i2;
    n7453_o2 <= n7453_i2;
    n7431_o2 <= n7431_i2;
    n7432_o2 <= n7432_i2;
    n7433_o2 <= n7433_i2;
    n7430_o2 <= n7430_i2;
    n7485_o2 <= n7485_i2;
    n7486_o2 <= n7486_i2;
    G2508_o2 <= G2508_i2;
    G2486_o2 <= G2486_i2;
    n2326_inv <= n7245_i2;
    n2329_inv <= n7246_i2;
    n3756_lo_buf_o2 <= n3756_lo_buf_i2;
    n4056_lo_buf_o2 <= n4056_lo_buf_i2;
    G3474_o2 <= G3474_i2;
    n2341_inv <= G2817_i2;
    n7396_o2 <= n7396_i2;
    n7398_o2 <= n7398_i2;
    n7400_o2 <= n7400_i2;
    n7401_o2 <= n7401_i2;
    n7402_o2 <= n7402_i2;
    n7403_o2 <= n7403_i2;
    n7404_o2 <= n7404_i2;
    n7405_o2 <= n7405_i2;
    G2711_o2 <= G2711_i2;
    n2371_inv <= G2828_i2;
    n7490_o2 <= n7490_i2;
    n7527_o2 <= n7527_i2;
    n7528_o2 <= n7528_i2;
    n7529_o2 <= n7529_i2;
    n7530_o2 <= n7530_i2;
    n7523_o2 <= n7523_i2;
    n7524_o2 <= n7524_i2;
    n7525_o2 <= n7525_i2;
    n7526_o2 <= n7526_i2;
    n4296_lo_buf_o2 <= n4296_lo_buf_i2;
    n4368_lo_buf_o2 <= n4368_lo_buf_i2;
    G2466_o2 <= G2466_i2;
    G2404_o2 <= G2404_i2;
    n7534_o2 <= n7534_i2;
    n7535_o2 <= n7535_i2;
    n7536_o2 <= n7536_i2;
    n7533_o2 <= n7533_i2;
    G1060_o2 <= G1060_i2;
    G963_o2 <= G963_i2;
    G2448_o2 <= G2448_i2;
    G2685_o2 <= G2685_i2;
    G2679_o2 <= G2679_i2;
    G2774_o2 <= G2774_i2;
    G2780_o2 <= G2780_i2;
    G2759_o2 <= G2759_i2;
    G2737_o2 <= G2737_i2;
    G2850_o2 <= G2850_i2;
    G3393_o2 <= G3393_i2;
    G3404_o2 <= G3404_i2;
    G3559_o2 <= G3559_i2;
    G2744_o2 <= G2744_i2;
    n3708_lo_buf_o2 <= n3708_lo_buf_i2;
    n3840_lo_buf_o2 <= n3840_lo_buf_i2;
    n4008_lo_buf_o2 <= n4008_lo_buf_i2;
    n4104_lo_buf_o2 <= n4104_lo_buf_i2;
    G1821_o2 <= G1821_i2;
    G1734_o2 <= G1734_i2;
    G3517_o2 <= G3517_i2;
    G3533_o2 <= G3533_i2;
    G3629_o2 <= G3629_i2;
    G3645_o2 <= G3645_i2;
    n2497_inv <= G2857_i2;
    G2731_o2 <= G2731_i2;
    G2844_o2 <= G2844_i2;
    n3732_lo_buf_o2 <= n3732_lo_buf_i2;
    n4032_lo_buf_o2 <= n4032_lo_buf_i2;
    G3552_o2 <= G3552_i2;
    G2271_o2 <= G2271_i2;
    n4248_lo_buf_o2 <= n4248_lo_buf_i2;
    n4332_lo_buf_o2 <= n4332_lo_buf_i2;
    n4344_lo_buf_o2 <= n4344_lo_buf_i2;
    n4380_lo_buf_o2 <= n4380_lo_buf_i2;
    G2398_o2 <= G2398_i2;
    G2480_o2 <= G2480_i2;
    G2418_o2 <= G2418_i2;
    G1455_o2 <= G1455_i2;
    G1449_o2 <= G1449_i2;
    G1452_o2 <= G1452_i2;
    G1425_o2 <= G1425_i2;
    G1428_o2 <= G1428_i2;
    G1419_o2 <= G1419_i2;
    G1422_o2 <= G1422_i2;
    n4308_lo_buf_o2 <= n4308_lo_buf_i2;
    G2675_o2 <= G2675_i2;
    G3035_o2 <= G3035_i2;
    G3026_o2 <= G3026_i2;
    G3029_o2 <= G3029_i2;
    G3032_o2 <= G3032_i2;
    G2999_o2 <= G2999_i2;
    G3002_o2 <= G3002_i2;
    G2770_o2 <= G2770_i2;
    G3008_o2 <= G3008_i2;
    G2073_o2 <= G2073_i2;
    G2752_o2 <= G2752_i2;
    G3005_o2 <= G3005_i2;
    G5108_o2 <= G5108_i2;
    G5135_o2 <= G5135_i2;
    G5111_o2 <= G5111_i2;
    G5138_o2 <= G5138_i2;
    G3415_o2 <= G3415_i2;
    G3386_o2 <= G3386_i2;
    G3570_o2 <= G3570_i2;
    G2430_o2 <= G2430_i2;
    G3495_o2 <= G3495_i2;
    G3621_o2 <= G3621_i2;
    n4284_lo_buf_o2 <= n4284_lo_buf_i2;
    n4356_lo_buf_o2 <= n4356_lo_buf_i2;
    G2472_o2 <= G2472_i2;
    G2410_o2 <= G2410_i2;
    n3960_lo_buf_o2 <= n3960_lo_buf_i2;
    n3972_lo_buf_o2 <= n3972_lo_buf_i2;
    n2647_inv <= G2865_i2;
    n2650_inv <= G970_i2;
    n3684_lo_buf_o2 <= n3684_lo_buf_i2;
    n4080_lo_buf_o2 <= n4080_lo_buf_i2;
    n4092_lo_buf_o2 <= n4092_lo_buf_i2;
    n2662_inv <= G1053_i2;
    n2665_inv <= G956_i2;
    G1147_o2 <= G1147_i2;
    G2705_o2 <= G2705_i2;
    G2693_o2 <= G2693_i2;
    G2696_o2 <= G2696_i2;
    G2700_o2 <= G2700_i2;
    G2915_o2 <= G2915_i2;
    G2966_o2 <= G2966_i2;
    G2540_o2 <= G2540_i2;
    G2788_o2 <= G2788_i2;
    G2792_o2 <= G2792_i2;
    G2797_o2 <= G2797_i2;
    G2804_o2 <= G2804_i2;
    G1038_o2 <= G1038_i2;
    G1044_o2 <= G1044_i2;
    G1090_o2 <= G1090_i2;
    G1096_o2 <= G1096_i2;
    G1029_o2 <= G1029_i2;
    G3942_o2 <= G3942_i2;
    G3954_o2 <= G3954_i2;
    G4011_o2 <= G4011_i2;
    G4017_o2 <= G4017_i2;
    G1141_o2 <= G1141_i2;
    G1081_o2 <= G1081_i2;
    G2146_o2 <= G2146_i2;
    G2145_o2 <= G2145_i2;
    G2144_o2 <= G2144_i2;
    G2143_o2 <= G2143_i2;
    G2142_o2 <= G2142_i2;
    G2141_o2 <= G2141_i2;
    G2140_o2 <= G2140_i2;
    G2139_o2 <= G2139_i2;
    G3769_o2 <= G3769_i2;
    G3773_o2 <= G3773_i2;
    G3768_o2 <= G3768_i2;
    G4101_o2 <= G4101_i2;
    G3161_o2 <= G3161_i2;
    G4143_o2 <= G4143_i2;
    G3828_o2 <= G3828_i2;
    G3831_o2 <= G3831_i2;
    G3334_o2 <= G3334_i2;
    G3335_o2 <= G3335_i2;
    G3180_o2 <= G3180_i2;
    G3340_o2 <= G3340_i2;
    G3339_o2 <= G3339_i2;
    G3341_o2 <= G3341_i2;
    G3234_o2 <= G3234_i2;
    G3829_o2 <= G3829_i2;
    G3338_o2 <= G3338_i2;
    G3336_o2 <= G3336_i2;
    G3770_o2 <= G3770_i2;
    G3918_o2 <= G3918_i2;
    G3774_o2 <= G3774_i2;
    G3921_o2 <= G3921_i2;
    G3832_o2 <= G3832_i2;
    G3993_o2 <= G3993_i2;
    G2076_o2 <= G2076_i2;
    G2071_o2 <= G2071_i2;
    G2072_o2 <= G2072_i2;
    G2069_o2 <= G2069_i2;
    G2070_o2 <= G2070_i2;
    G2067_o2 <= G2067_i2;
    G2068_o2 <= G2068_i2;
    G4095_o2 <= G4095_i2;
    G3272_o2 <= G3272_i2;
    G3269_o2 <= G3269_i2;
    G3270_o2 <= G3270_i2;
    G3271_o2 <= G3271_i2;
    G3265_o2 <= G3265_i2;
    G3266_o2 <= G3266_i2;
    G4137_o2 <= G4137_i2;
    G3268_o2 <= G3268_i2;
    G2361_o2 <= G2361_i2;
    G3228_o2 <= G3228_i2;
    G3267_o2 <= G3267_i2;
    G2336_o2 <= G2336_i2;
    G3459_o2 <= G3459_i2;
    G3428_o2 <= G3428_i2;
    G3438_o2 <= G3438_i2;
    G3449_o2 <= G3449_i2;
    G3421_o2 <= G3421_i2;
    G3576_o2 <= G3576_i2;
    G3303_o2 <= G3303_i2;
    G3583_o2 <= G3583_i2;
    G3594_o2 <= G3594_i2;
    G3674_o2 <= G3674_i2;
    G3685_o2 <= G3685_i2;
    G4504_o2 <= G4504_i2;
    G4180_o2 <= G4180_i2;
    G5123_o2 <= G5123_i2;
    G5142_o2 <= G5142_i2;
    G5126_o2 <= G5126_i2;
    G5144_o2 <= G5144_i2;
    G3912_o2 <= G3912_i2;
    G4417_o2 <= G4417_i2;
    G4420_o2 <= G4420_i2;
    G3969_o2 <= G3969_i2;
    G4023_o2 <= G4023_i2;
    G2720_o2 <= G2720_i2;
    G2837_o2 <= G2837_i2;
    n2965_inv <= G836_i2;
    n2968_inv <= G848_i2;
    n2971_inv <= G813_i2;
    n2974_inv <= G825_i2;
    G1876_o2 <= G1876_i2;
    G4996_o2 <= G4996_i2;
    G4984_o2 <= G4984_i2;
    G4920_o2 <= G4920_i2;
    G4923_o2 <= G4923_i2;
    G4930_o2 <= G4930_i2;
    G4933_o2 <= G4933_i2;
    n4320_lo_buf_o2 <= n4320_lo_buf_i2;
    G2424_o2 <= G2424_i2;
    G3317_o2 <= G3317_i2;
    G3503_o2 <= G3503_i2;
    G3485_o2 <= G3485_i2;
    G3611_o2 <= G3611_i2;
    n3864_lo_buf_o2 <= n3864_lo_buf_i2;
    n3888_lo_buf_o2 <= n3888_lo_buf_i2;
    n4116_lo_buf_o2 <= n4116_lo_buf_i2;
    n4128_lo_buf_o2 <= n4128_lo_buf_i2;
    n4140_lo_buf_o2 <= n4140_lo_buf_i2;
    n4152_lo_buf_o2 <= n4152_lo_buf_i2;
    G1815_o2 <= G1815_i2;
    G1728_o2 <= G1728_i2;
    G1035_o2 <= G1035_i2;
    G1041_o2 <= G1041_i2;
    G1087_o2 <= G1087_i2;
    G1093_o2 <= G1093_i2;
    G1132_o2 <= G1132_i2;
    G1108_o2 <= G1108_i2;
    G1138_o2 <= G1138_i2;
    G1114_o2 <= G1114_i2;
    G1807_o2 <= G1807_i2;
    G2108_o2 <= G2108_i2;
    G1126_o2 <= G1126_i2;
    G1899_o2 <= G1899_i2;
    G2134_o2 <= G2134_i2;
    G1852_o2 <= G1852_i2;
    G2116_o2 <= G2116_i2;
    G2543_o2 <= G2543_i2;
    G2727_o2 <= G2727_i2;
    G2715_o2 <= G2715_i2;
    G2832_o2 <= G2832_i2;
    G1873_o2 <= G1873_i2;
    G3291_o2 <= G3291_i2;
    G5025_o2 <= G5025_i2;
    G5036_o2 <= G5036_i2;
    G3132_o2 <= G3132_i2;
    G5038_o2 <= G5038_i2;
    G5039_o2 <= G5039_i2;
    n3118_inv <= G1150_i2;
    n3121_inv <= G1162_i2;
    n3124_inv <= G804_i2;
    n3127_inv <= G1172_i2;
    n3984_lo_buf_o2 <= n3984_lo_buf_i2;
    G1802_o2 <= G1802_i2;
    G1804_o2 <= G1804_i2;
    G1849_o2 <= G1849_i2;
    G1851_o2 <= G1851_i2;
    G2492_o2 <= G2492_i2;
    G1799_o2 <= G1799_i2;
    G4231_o2 <= G4231_i2;
    G4234_o2 <= G4234_i2;
    G4245_o2 <= G4245_i2;
    G4247_o2 <= G4247_i2;
    G1894_o2 <= G1894_i2;
    G1846_o2 <= G1846_i2;
    G4238_o2 <= G4238_i2;
    G4249_o2 <= G4249_i2;
    G2293_o2 <= G2293_i2;
    G5022_o2 <= G5022_i2;
    G5006_o2 <= G5006_i2;
    G4944_o2 <= G4944_i2;
    G4946_o2 <= G4946_i2;
    G4954_o2 <= G4954_i2;
    G4956_o2 <= G4956_i2;
    G3546_o2 <= G3546_i2;
    G3658_o2 <= G3658_i2;
    G1344_o2 <= G1344_i2;
    G2921_o2 <= G2921_i2;
    n3912_lo_buf_o2 <= n3912_lo_buf_i2;
    G1835_o2 <= G1835_i2;
    G3810_o2 <= G3810_i2;
    G3866_o2 <= G3866_i2;
    G3811_o2 <= G3811_i2;
    G2269_o2 <= G2269_i2;
    G3812_o2 <= G3812_i2;
    G3867_o2 <= G3867_i2;
    G3868_o2 <= G3868_i2;
    G3809_o2 <= G3809_i2;
    G3716_o2 <= G3716_i2;
    G4529_o2 <= G4529_i2;
    G4670_o2 <= G4670_i2;
    G4493_o2 <= G4493_i2;
    G4580_o2 <= G4580_i2;
    G3822_o2 <= G3822_i2;
    G3877_o2 <= G3877_i2;
    G4131_o2 <= G4131_i2;
    G4170_o2 <= G4170_i2;
    G4051_o2 <= G4051_i2;
    G4065_o2 <= G4065_i2;
    G4697_o2 <= G4697_i2;
    G4706_o2 <= G4706_i2;
    G2460_o2 <= G2460_i2;
    G2454_o2 <= G2454_i2;
    G2392_o2 <= G2392_i2;
    G2386_o2 <= G2386_i2;
    n4260_lo_buf_o2 <= n4260_lo_buf_i2;
    n4272_lo_buf_o2 <= n4272_lo_buf_i2;
    n4392_lo_buf_o2 <= n4392_lo_buf_i2;
    n4404_lo_buf_o2 <= n4404_lo_buf_i2;
    G1512_o2 <= G1512_i2;
    G3135_o2 <= G3135_i2;
    G2379_o2 <= G2379_i2;
    n4164_lo_buf_o2 <= n4164_lo_buf_i2;
    n4176_lo_buf_o2 <= n4176_lo_buf_i2;
    n4224_lo_buf_o2 <= n4224_lo_buf_i2;
    G2975_o2 <= G2975_i2;
    G2978_o2 <= G2978_i2;
    G2933_o2 <= G2933_i2;
    G2936_o2 <= G2936_i2;
    G1356_o2 <= G1356_i2;
    G1359_o2 <= G1359_i2;
    G1398_o2 <= G1398_i2;
    G1401_o2 <= G1401_i2;
  end
  initial begin
    n2610_lo <= 1'b0;
    n2613_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2622_lo <= 1'b0;
    n2625_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2631_lo <= 1'b0;
    n2634_lo <= 1'b0;
    n2637_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2646_lo <= 1'b0;
    n2649_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2658_lo <= 1'b0;
    n2661_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2670_lo <= 1'b0;
    n2673_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2694_lo <= 1'b0;
    n2697_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2706_lo <= 1'b0;
    n2709_lo <= 1'b0;
    n2712_lo <= 1'b0;
    n2715_lo <= 1'b0;
    n2718_lo <= 1'b0;
    n2721_lo <= 1'b0;
    n2724_lo <= 1'b0;
    n2727_lo <= 1'b0;
    n2730_lo <= 1'b0;
    n2733_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2742_lo <= 1'b0;
    n2745_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2754_lo <= 1'b0;
    n2757_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2766_lo <= 1'b0;
    n2769_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2778_lo <= 1'b0;
    n2781_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2811_lo <= 1'b0;
    n2814_lo <= 1'b0;
    n2817_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2847_lo <= 1'b0;
    n2850_lo <= 1'b0;
    n2853_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2910_lo <= 1'b0;
    n2913_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2922_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2931_lo <= 1'b0;
    n2934_lo <= 1'b0;
    n2937_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2946_lo <= 1'b0;
    n2949_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2958_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2973_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2985_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3009_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3042_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3066_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3078_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3090_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3144_lo <= 1'b0;
    n3147_lo <= 1'b0;
    n3150_lo <= 1'b0;
    n3153_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3159_lo <= 1'b0;
    n3162_lo <= 1'b0;
    n3165_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3186_lo <= 1'b0;
    n3189_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3198_lo <= 1'b0;
    n3201_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3213_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3225_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3234_lo <= 1'b0;
    n3237_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3246_lo <= 1'b0;
    n3249_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3261_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3273_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3285_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3297_lo <= 1'b0;
    n3300_lo <= 1'b0;
    n3303_lo <= 1'b0;
    n3306_lo <= 1'b0;
    n3309_lo <= 1'b0;
    n3312_lo <= 1'b0;
    n3315_lo <= 1'b0;
    n3318_lo <= 1'b0;
    n3321_lo <= 1'b0;
    n3324_lo <= 1'b0;
    n3327_lo <= 1'b0;
    n3330_lo <= 1'b0;
    n3333_lo <= 1'b0;
    n3336_lo <= 1'b0;
    n3339_lo <= 1'b0;
    n3342_lo <= 1'b0;
    n3345_lo <= 1'b0;
    n3348_lo <= 1'b0;
    n3351_lo <= 1'b0;
    n3354_lo <= 1'b0;
    n3357_lo <= 1'b0;
    n3360_lo <= 1'b0;
    n3363_lo <= 1'b0;
    n3366_lo <= 1'b0;
    n3369_lo <= 1'b0;
    n3372_lo <= 1'b0;
    n3375_lo <= 1'b0;
    n3378_lo <= 1'b0;
    n3381_lo <= 1'b0;
    n3384_lo <= 1'b0;
    n3387_lo <= 1'b0;
    n3390_lo <= 1'b0;
    n3393_lo <= 1'b0;
    n3396_lo <= 1'b0;
    n3399_lo <= 1'b0;
    n3402_lo <= 1'b0;
    n3405_lo <= 1'b0;
    n3408_lo <= 1'b0;
    n3411_lo <= 1'b0;
    n3414_lo <= 1'b0;
    n3417_lo <= 1'b0;
    n3420_lo <= 1'b0;
    n3423_lo <= 1'b0;
    n3426_lo <= 1'b0;
    n3429_lo <= 1'b0;
    n3432_lo <= 1'b0;
    n3435_lo <= 1'b0;
    n3438_lo <= 1'b0;
    n3441_lo <= 1'b0;
    n3444_lo <= 1'b0;
    n3447_lo <= 1'b0;
    n3450_lo <= 1'b0;
    n3453_lo <= 1'b0;
    n3456_lo <= 1'b0;
    n3459_lo <= 1'b0;
    n3462_lo <= 1'b0;
    n3465_lo <= 1'b0;
    n3468_lo <= 1'b0;
    n3471_lo <= 1'b0;
    n3474_lo <= 1'b0;
    n3477_lo <= 1'b0;
    n3480_lo <= 1'b0;
    n3483_lo <= 1'b0;
    n3486_lo <= 1'b0;
    n3489_lo <= 1'b0;
    n3492_lo <= 1'b0;
    n3495_lo <= 1'b0;
    n3498_lo <= 1'b0;
    n3501_lo <= 1'b0;
    n3504_lo <= 1'b0;
    n3507_lo <= 1'b0;
    n3510_lo <= 1'b0;
    n3513_lo <= 1'b0;
    n3516_lo <= 1'b0;
    n3519_lo <= 1'b0;
    n3522_lo <= 1'b0;
    n3525_lo <= 1'b0;
    n3528_lo <= 1'b0;
    n3531_lo <= 1'b0;
    n3534_lo <= 1'b0;
    n3537_lo <= 1'b0;
    n3540_lo <= 1'b0;
    n3543_lo <= 1'b0;
    n3546_lo <= 1'b0;
    n3549_lo <= 1'b0;
    n3552_lo <= 1'b0;
    n3555_lo <= 1'b0;
    n3558_lo <= 1'b0;
    n3561_lo <= 1'b0;
    n3564_lo <= 1'b0;
    n3567_lo <= 1'b0;
    n3570_lo <= 1'b0;
    n3573_lo <= 1'b0;
    n3576_lo <= 1'b0;
    n3579_lo <= 1'b0;
    n3582_lo <= 1'b0;
    n3585_lo <= 1'b0;
    n3588_lo <= 1'b0;
    n3591_lo <= 1'b0;
    n3594_lo <= 1'b0;
    n3597_lo <= 1'b0;
    n3600_lo <= 1'b0;
    n3603_lo <= 1'b0;
    n3606_lo <= 1'b0;
    n3609_lo <= 1'b0;
    n3612_lo <= 1'b0;
    n3615_lo <= 1'b0;
    n3618_lo <= 1'b0;
    n3621_lo <= 1'b0;
    n3624_lo <= 1'b0;
    n3627_lo <= 1'b0;
    n3630_lo <= 1'b0;
    n3633_lo <= 1'b0;
    n3636_lo <= 1'b0;
    n3639_lo <= 1'b0;
    n3642_lo <= 1'b0;
    n3645_lo <= 1'b0;
    n3648_lo <= 1'b0;
    n3651_lo <= 1'b0;
    n3654_lo <= 1'b0;
    n3657_lo <= 1'b0;
    n3666_lo <= 1'b0;
    n3669_lo <= 1'b0;
    n3678_lo <= 1'b0;
    n3687_lo <= 1'b0;
    n3690_lo <= 1'b0;
    n3702_lo <= 1'b0;
    n3711_lo <= 1'b0;
    n3714_lo <= 1'b0;
    n3726_lo <= 1'b0;
    n3735_lo <= 1'b0;
    n3738_lo <= 1'b0;
    n3750_lo <= 1'b0;
    n3753_lo <= 1'b0;
    n3759_lo <= 1'b0;
    n3762_lo <= 1'b0;
    n3765_lo <= 1'b0;
    n3774_lo <= 1'b0;
    n3777_lo <= 1'b0;
    n3786_lo <= 1'b0;
    n3789_lo <= 1'b0;
    n3792_lo <= 1'b0;
    n3795_lo <= 1'b0;
    n3798_lo <= 1'b0;
    n3801_lo <= 1'b0;
    n3810_lo <= 1'b0;
    n3813_lo <= 1'b0;
    n3822_lo <= 1'b0;
    n3825_lo <= 1'b0;
    n3834_lo <= 1'b0;
    n3843_lo <= 1'b0;
    n3846_lo <= 1'b0;
    n3867_lo <= 1'b0;
    n3891_lo <= 1'b0;
    n3915_lo <= 1'b0;
    n3930_lo <= 1'b0;
    n3933_lo <= 1'b0;
    n3936_lo <= 1'b0;
    n3942_lo <= 1'b0;
    n3945_lo <= 1'b0;
    n3948_lo <= 1'b0;
    n3954_lo <= 1'b0;
    n3957_lo <= 1'b0;
    n3963_lo <= 1'b0;
    n3966_lo <= 1'b0;
    n3969_lo <= 1'b0;
    n3975_lo <= 1'b0;
    n3978_lo <= 1'b0;
    n3987_lo <= 1'b0;
    n3990_lo <= 1'b0;
    n4002_lo <= 1'b0;
    n4011_lo <= 1'b0;
    n4014_lo <= 1'b0;
    n4026_lo <= 1'b0;
    n4035_lo <= 1'b0;
    n4038_lo <= 1'b0;
    n4050_lo <= 1'b0;
    n4053_lo <= 1'b0;
    n4059_lo <= 1'b0;
    n4062_lo <= 1'b0;
    n4065_lo <= 1'b0;
    n4098_lo <= 1'b0;
    n4107_lo <= 1'b0;
    n4119_lo <= 1'b0;
    n4131_lo <= 1'b0;
    n4143_lo <= 1'b0;
    n4155_lo <= 1'b0;
    n4167_lo <= 1'b0;
    n4179_lo <= 1'b0;
    n4182_lo <= 1'b0;
    n4185_lo <= 1'b0;
    n4188_lo <= 1'b0;
    n4194_lo <= 1'b0;
    n4197_lo <= 1'b0;
    n4200_lo <= 1'b0;
    n4206_lo <= 1'b0;
    n4209_lo <= 1'b0;
    n4212_lo <= 1'b0;
    n4215_lo <= 1'b0;
    n4227_lo <= 1'b0;
    n4230_lo <= 1'b0;
    n4233_lo <= 1'b0;
    n4236_lo <= 1'b0;
    n4239_lo <= 1'b0;
    n4242_lo <= 1'b0;
    n4251_lo <= 1'b0;
    n4263_lo <= 1'b0;
    n4275_lo <= 1'b0;
    n4278_lo <= 1'b0;
    n4287_lo <= 1'b0;
    n4290_lo <= 1'b0;
    n4293_lo <= 1'b0;
    n4299_lo <= 1'b0;
    n4302_lo <= 1'b0;
    n4305_lo <= 1'b0;
    n4311_lo <= 1'b0;
    n4314_lo <= 1'b0;
    n4323_lo <= 1'b0;
    n4326_lo <= 1'b0;
    n4335_lo <= 1'b0;
    n4338_lo <= 1'b0;
    n4347_lo <= 1'b0;
    n4350_lo <= 1'b0;
    n4359_lo <= 1'b0;
    n4362_lo <= 1'b0;
    n4365_lo <= 1'b0;
    n4371_lo <= 1'b0;
    n4374_lo <= 1'b0;
    n4383_lo <= 1'b0;
    n4395_lo <= 1'b0;
    n4407_lo <= 1'b0;
    n4410_lo <= 1'b0;
    n4413_lo <= 1'b0;
    n4416_lo <= 1'b0;
    n4419_lo <= 1'b0;
    n4422_lo <= 1'b0;
    n4425_lo <= 1'b0;
    n4428_lo <= 1'b0;
    n4431_lo <= 1'b0;
    n4434_lo <= 1'b0;
    n4437_lo <= 1'b0;
    n4440_lo <= 1'b0;
    n4443_lo <= 1'b0;
    n4446_lo <= 1'b0;
    n4449_lo <= 1'b0;
    n4452_lo <= 1'b0;
    n4455_lo <= 1'b0;
    n4458_lo <= 1'b0;
    n4461_lo <= 1'b0;
    n4464_lo <= 1'b0;
    n4467_lo <= 1'b0;
    n4470_lo <= 1'b0;
    n4473_lo <= 1'b0;
    n4476_lo <= 1'b0;
    n4479_lo <= 1'b0;
    n4482_lo <= 1'b0;
    n4485_lo <= 1'b0;
    n4488_lo <= 1'b0;
    n4494_lo <= 1'b0;
    n4497_lo <= 1'b0;
    n4500_lo <= 1'b0;
    n4503_lo <= 1'b0;
    n4506_lo <= 1'b0;
    n4509_lo <= 1'b0;
    n4512_lo <= 1'b0;
    n4515_lo <= 1'b0;
    n4518_lo <= 1'b0;
    n4521_lo <= 1'b0;
    n4524_lo <= 1'b0;
    n4527_lo <= 1'b0;
    n4530_lo <= 1'b0;
    n4533_lo <= 1'b0;
    n4536_lo <= 1'b0;
    n4539_lo <= 1'b0;
    n4542_lo <= 1'b0;
    n4545_lo <= 1'b0;
    n4548_lo <= 1'b0;
    n4554_lo <= 1'b0;
    n4557_lo <= 1'b0;
    n4560_lo <= 1'b0;
    n4563_lo <= 1'b0;
    n4566_lo <= 1'b0;
    n4569_lo <= 1'b0;
    n4572_lo <= 1'b0;
    n4575_lo <= 1'b0;
    n4578_lo <= 1'b0;
    n4581_lo <= 1'b0;
    n4584_lo <= 1'b0;
    n4587_lo <= 1'b0;
    n4590_lo <= 1'b0;
    n4593_lo <= 1'b0;
    n4596_lo <= 1'b0;
    n4599_lo <= 1'b0;
    n4602_lo <= 1'b0;
    n4605_lo <= 1'b0;
    n4608_lo <= 1'b0;
    n4611_lo <= 1'b0;
    n4614_lo <= 1'b0;
    n4617_lo <= 1'b0;
    n4620_lo <= 1'b0;
    n4623_lo <= 1'b0;
    n4626_lo <= 1'b0;
    n4629_lo <= 1'b0;
    n4632_lo <= 1'b0;
    n4635_lo <= 1'b0;
    n4638_lo <= 1'b0;
    n4641_lo <= 1'b0;
    n4644_lo <= 1'b0;
    n4647_lo <= 1'b0;
    n4650_lo <= 1'b0;
    n4653_lo <= 1'b0;
    n4656_lo <= 1'b0;
    n4659_lo <= 1'b0;
    n4662_lo <= 1'b0;
    n4665_lo <= 1'b0;
    n4668_lo <= 1'b0;
    n4671_lo <= 1'b0;
    n4674_lo <= 1'b0;
    n4677_lo <= 1'b0;
    n4680_lo <= 1'b0;
    n4683_lo <= 1'b0;
    n4686_lo <= 1'b0;
    n4689_lo <= 1'b0;
    n4692_lo <= 1'b0;
    n4695_lo <= 1'b0;
    n4698_lo <= 1'b0;
    n4701_lo <= 1'b0;
    n4704_lo <= 1'b0;
    n4707_lo <= 1'b0;
    n4710_lo <= 1'b0;
    n4713_lo <= 1'b0;
    n4716_lo <= 1'b0;
    n4719_lo <= 1'b0;
    n4722_lo <= 1'b0;
    n4725_lo <= 1'b0;
    n4728_lo <= 1'b0;
    n4731_lo <= 1'b0;
    n4734_lo <= 1'b0;
    n4737_lo <= 1'b0;
    n4740_lo <= 1'b0;
    n4743_lo <= 1'b0;
    n6382_o2 <= 1'b0;
    n6383_o2 <= 1'b0;
    n6419_o2 <= 1'b0;
    n6420_o2 <= 1'b0;
    n6435_o2 <= 1'b0;
    n6436_o2 <= 1'b0;
    n6448_o2 <= 1'b0;
    n6449_o2 <= 1'b0;
    n6613_o2 <= 1'b0;
    n6614_o2 <= 1'b0;
    n6641_o2 <= 1'b0;
    n6658_o2 <= 1'b0;
    n6757_o2 <= 1'b0;
    n6756_o2 <= 1'b0;
    n7116_o2 <= 1'b0;
    n7156_o2 <= 1'b0;
    n6549_o2 <= 1'b0;
    n6550_o2 <= 1'b0;
    n7357_o2 <= 1'b0;
    n7358_o2 <= 1'b0;
    n7359_o2 <= 1'b0;
    n7360_o2 <= 1'b0;
    n6621_o2 <= 1'b0;
    n6623_o2 <= 1'b0;
    n6625_o2 <= 1'b0;
    n6626_o2 <= 1'b0;
    n6627_o2 <= 1'b0;
    n6628_o2 <= 1'b0;
    n6629_o2 <= 1'b0;
    n6630_o2 <= 1'b0;
    n6669_o2 <= 1'b0;
    n7449_o2 <= 1'b0;
    n7450_o2 <= 1'b0;
    n7451_o2 <= 1'b0;
    n7452_o2 <= 1'b0;
    n6682_o2 <= 1'b0;
    n6683_o2 <= 1'b0;
    n6684_o2 <= 1'b0;
    n6685_o2 <= 1'b0;
    n7463_o2 <= 1'b0;
    n6686_o2 <= 1'b0;
    n6687_o2 <= 1'b0;
    n6688_o2 <= 1'b0;
    n6689_o2 <= 1'b0;
    n6772_o2 <= 1'b0;
    n6773_o2 <= 1'b0;
    n6774_o2 <= 1'b0;
    n6775_o2 <= 1'b0;
    G3467_o2 <= 1'b0;
    G2810_o2 <= 1'b0;
    n6833_o2 <= 1'b0;
    n6945_o2 <= 1'b0;
    n6947_o2 <= 1'b0;
    n6949_o2 <= 1'b0;
    n6951_o2 <= 1'b0;
    n6888_o2 <= 1'b0;
    n6889_o2 <= 1'b0;
    n6936_o2 <= 1'b0;
    n6954_o2 <= 1'b0;
    n6955_o2 <= 1'b0;
    n6956_o2 <= 1'b0;
    n6957_o2 <= 1'b0;
    n6958_o2 <= 1'b0;
    n6982_o2 <= 1'b0;
    n6984_o2 <= 1'b0;
    n6974_o2 <= 1'b0;
    n6975_o2 <= 1'b0;
    n6999_o2 <= 1'b0;
    n7015_o2 <= 1'b0;
    n7016_o2 <= 1'b0;
    n7017_o2 <= 1'b0;
    n7018_o2 <= 1'b0;
    n7005_o2 <= 1'b0;
    n7019_o2 <= 1'b0;
    n7022_o2 <= 1'b0;
    n7023_o2 <= 1'b0;
    n7132_o2 <= 1'b0;
    n7133_o2 <= 1'b0;
    n7135_o2 <= 1'b0;
    n7136_o2 <= 1'b0;
    n7175_o2 <= 1'b0;
    n7155_o2 <= 1'b0;
    G3060_o2 <= 1'b0;
    n7383_o2 <= 1'b0;
    G3802_o2 <= 1'b0;
    G3859_o2 <= 1'b0;
    n7355_o2 <= 1'b0;
    n7356_o2 <= 1'b0;
    G4054_o2 <= 1'b0;
    G4068_o2 <= 1'b0;
    n7384_o2 <= 1'b0;
    n7387_o2 <= 1'b0;
    n7388_o2 <= 1'b0;
    n7389_o2 <= 1'b0;
    n7386_o2 <= 1'b0;
    n7453_o2 <= 1'b0;
    n7431_o2 <= 1'b0;
    n7432_o2 <= 1'b0;
    n7433_o2 <= 1'b0;
    n7430_o2 <= 1'b0;
    n7485_o2 <= 1'b0;
    n7486_o2 <= 1'b0;
    G2508_o2 <= 1'b0;
    G2486_o2 <= 1'b0;
    n2326_inv <= 1'b0;
    n2329_inv <= 1'b0;
    n3756_lo_buf_o2 <= 1'b0;
    n4056_lo_buf_o2 <= 1'b0;
    G3474_o2 <= 1'b0;
    n2341_inv <= 1'b0;
    n7396_o2 <= 1'b0;
    n7398_o2 <= 1'b0;
    n7400_o2 <= 1'b0;
    n7401_o2 <= 1'b0;
    n7402_o2 <= 1'b0;
    n7403_o2 <= 1'b0;
    n7404_o2 <= 1'b0;
    n7405_o2 <= 1'b0;
    G2711_o2 <= 1'b0;
    n2371_inv <= 1'b0;
    n7490_o2 <= 1'b0;
    n7527_o2 <= 1'b0;
    n7528_o2 <= 1'b0;
    n7529_o2 <= 1'b0;
    n7530_o2 <= 1'b0;
    n7523_o2 <= 1'b0;
    n7524_o2 <= 1'b0;
    n7525_o2 <= 1'b0;
    n7526_o2 <= 1'b0;
    n4296_lo_buf_o2 <= 1'b0;
    n4368_lo_buf_o2 <= 1'b0;
    G2466_o2 <= 1'b0;
    G2404_o2 <= 1'b0;
    n7534_o2 <= 1'b0;
    n7535_o2 <= 1'b0;
    n7536_o2 <= 1'b0;
    n7533_o2 <= 1'b0;
    G1060_o2 <= 1'b0;
    G963_o2 <= 1'b0;
    G2448_o2 <= 1'b0;
    G2685_o2 <= 1'b0;
    G2679_o2 <= 1'b0;
    G2774_o2 <= 1'b0;
    G2780_o2 <= 1'b0;
    G2759_o2 <= 1'b0;
    G2737_o2 <= 1'b0;
    G2850_o2 <= 1'b0;
    G3393_o2 <= 1'b0;
    G3404_o2 <= 1'b0;
    G3559_o2 <= 1'b0;
    G2744_o2 <= 1'b0;
    n3708_lo_buf_o2 <= 1'b0;
    n3840_lo_buf_o2 <= 1'b0;
    n4008_lo_buf_o2 <= 1'b0;
    n4104_lo_buf_o2 <= 1'b0;
    G1821_o2 <= 1'b0;
    G1734_o2 <= 1'b0;
    G3517_o2 <= 1'b0;
    G3533_o2 <= 1'b0;
    G3629_o2 <= 1'b0;
    G3645_o2 <= 1'b0;
    n2497_inv <= 1'b0;
    G2731_o2 <= 1'b0;
    G2844_o2 <= 1'b0;
    n3732_lo_buf_o2 <= 1'b0;
    n4032_lo_buf_o2 <= 1'b0;
    G3552_o2 <= 1'b0;
    G2271_o2 <= 1'b0;
    n4248_lo_buf_o2 <= 1'b0;
    n4332_lo_buf_o2 <= 1'b0;
    n4344_lo_buf_o2 <= 1'b0;
    n4380_lo_buf_o2 <= 1'b0;
    G2398_o2 <= 1'b0;
    G2480_o2 <= 1'b0;
    G2418_o2 <= 1'b0;
    G1455_o2 <= 1'b0;
    G1449_o2 <= 1'b0;
    G1452_o2 <= 1'b0;
    G1425_o2 <= 1'b0;
    G1428_o2 <= 1'b0;
    G1419_o2 <= 1'b0;
    G1422_o2 <= 1'b0;
    n4308_lo_buf_o2 <= 1'b0;
    G2675_o2 <= 1'b0;
    G3035_o2 <= 1'b0;
    G3026_o2 <= 1'b0;
    G3029_o2 <= 1'b0;
    G3032_o2 <= 1'b0;
    G2999_o2 <= 1'b0;
    G3002_o2 <= 1'b0;
    G2770_o2 <= 1'b0;
    G3008_o2 <= 1'b0;
    G2073_o2 <= 1'b0;
    G2752_o2 <= 1'b0;
    G3005_o2 <= 1'b0;
    G5108_o2 <= 1'b0;
    G5135_o2 <= 1'b0;
    G5111_o2 <= 1'b0;
    G5138_o2 <= 1'b0;
    G3415_o2 <= 1'b0;
    G3386_o2 <= 1'b0;
    G3570_o2 <= 1'b0;
    G2430_o2 <= 1'b0;
    G3495_o2 <= 1'b0;
    G3621_o2 <= 1'b0;
    n4284_lo_buf_o2 <= 1'b0;
    n4356_lo_buf_o2 <= 1'b0;
    G2472_o2 <= 1'b0;
    G2410_o2 <= 1'b0;
    n3960_lo_buf_o2 <= 1'b0;
    n3972_lo_buf_o2 <= 1'b0;
    n2647_inv <= 1'b0;
    n2650_inv <= 1'b0;
    n3684_lo_buf_o2 <= 1'b0;
    n4080_lo_buf_o2 <= 1'b0;
    n4092_lo_buf_o2 <= 1'b0;
    n2662_inv <= 1'b0;
    n2665_inv <= 1'b0;
    G1147_o2 <= 1'b0;
    G2705_o2 <= 1'b0;
    G2693_o2 <= 1'b0;
    G2696_o2 <= 1'b0;
    G2700_o2 <= 1'b0;
    G2915_o2 <= 1'b0;
    G2966_o2 <= 1'b0;
    G2540_o2 <= 1'b0;
    G2788_o2 <= 1'b0;
    G2792_o2 <= 1'b0;
    G2797_o2 <= 1'b0;
    G2804_o2 <= 1'b0;
    G1038_o2 <= 1'b0;
    G1044_o2 <= 1'b0;
    G1090_o2 <= 1'b0;
    G1096_o2 <= 1'b0;
    G1029_o2 <= 1'b0;
    G3942_o2 <= 1'b0;
    G3954_o2 <= 1'b0;
    G4011_o2 <= 1'b0;
    G4017_o2 <= 1'b0;
    G1141_o2 <= 1'b0;
    G1081_o2 <= 1'b0;
    G2146_o2 <= 1'b0;
    G2145_o2 <= 1'b0;
    G2144_o2 <= 1'b0;
    G2143_o2 <= 1'b0;
    G2142_o2 <= 1'b0;
    G2141_o2 <= 1'b0;
    G2140_o2 <= 1'b0;
    G2139_o2 <= 1'b0;
    G3769_o2 <= 1'b0;
    G3773_o2 <= 1'b0;
    G3768_o2 <= 1'b0;
    G4101_o2 <= 1'b0;
    G3161_o2 <= 1'b0;
    G4143_o2 <= 1'b0;
    G3828_o2 <= 1'b0;
    G3831_o2 <= 1'b0;
    G3334_o2 <= 1'b0;
    G3335_o2 <= 1'b0;
    G3180_o2 <= 1'b0;
    G3340_o2 <= 1'b0;
    G3339_o2 <= 1'b0;
    G3341_o2 <= 1'b0;
    G3234_o2 <= 1'b0;
    G3829_o2 <= 1'b0;
    G3338_o2 <= 1'b0;
    G3336_o2 <= 1'b0;
    G3770_o2 <= 1'b0;
    G3918_o2 <= 1'b0;
    G3774_o2 <= 1'b0;
    G3921_o2 <= 1'b0;
    G3832_o2 <= 1'b0;
    G3993_o2 <= 1'b0;
    G2076_o2 <= 1'b0;
    G2071_o2 <= 1'b0;
    G2072_o2 <= 1'b0;
    G2069_o2 <= 1'b0;
    G2070_o2 <= 1'b0;
    G2067_o2 <= 1'b0;
    G2068_o2 <= 1'b0;
    G4095_o2 <= 1'b0;
    G3272_o2 <= 1'b0;
    G3269_o2 <= 1'b0;
    G3270_o2 <= 1'b0;
    G3271_o2 <= 1'b0;
    G3265_o2 <= 1'b0;
    G3266_o2 <= 1'b0;
    G4137_o2 <= 1'b0;
    G3268_o2 <= 1'b0;
    G2361_o2 <= 1'b0;
    G3228_o2 <= 1'b0;
    G3267_o2 <= 1'b0;
    G2336_o2 <= 1'b0;
    G3459_o2 <= 1'b0;
    G3428_o2 <= 1'b0;
    G3438_o2 <= 1'b0;
    G3449_o2 <= 1'b0;
    G3421_o2 <= 1'b0;
    G3576_o2 <= 1'b0;
    G3303_o2 <= 1'b0;
    G3583_o2 <= 1'b0;
    G3594_o2 <= 1'b0;
    G3674_o2 <= 1'b0;
    G3685_o2 <= 1'b0;
    G4504_o2 <= 1'b0;
    G4180_o2 <= 1'b0;
    G5123_o2 <= 1'b0;
    G5142_o2 <= 1'b0;
    G5126_o2 <= 1'b0;
    G5144_o2 <= 1'b0;
    G3912_o2 <= 1'b0;
    G4417_o2 <= 1'b0;
    G4420_o2 <= 1'b0;
    G3969_o2 <= 1'b0;
    G4023_o2 <= 1'b0;
    G2720_o2 <= 1'b0;
    G2837_o2 <= 1'b0;
    n2965_inv <= 1'b0;
    n2968_inv <= 1'b0;
    n2971_inv <= 1'b0;
    n2974_inv <= 1'b0;
    G1876_o2 <= 1'b0;
    G4996_o2 <= 1'b0;
    G4984_o2 <= 1'b0;
    G4920_o2 <= 1'b0;
    G4923_o2 <= 1'b0;
    G4930_o2 <= 1'b0;
    G4933_o2 <= 1'b0;
    n4320_lo_buf_o2 <= 1'b0;
    G2424_o2 <= 1'b0;
    G3317_o2 <= 1'b0;
    G3503_o2 <= 1'b0;
    G3485_o2 <= 1'b0;
    G3611_o2 <= 1'b0;
    n3864_lo_buf_o2 <= 1'b0;
    n3888_lo_buf_o2 <= 1'b0;
    n4116_lo_buf_o2 <= 1'b0;
    n4128_lo_buf_o2 <= 1'b0;
    n4140_lo_buf_o2 <= 1'b0;
    n4152_lo_buf_o2 <= 1'b0;
    G1815_o2 <= 1'b0;
    G1728_o2 <= 1'b0;
    G1035_o2 <= 1'b0;
    G1041_o2 <= 1'b0;
    G1087_o2 <= 1'b0;
    G1093_o2 <= 1'b0;
    G1132_o2 <= 1'b0;
    G1108_o2 <= 1'b0;
    G1138_o2 <= 1'b0;
    G1114_o2 <= 1'b0;
    G1807_o2 <= 1'b0;
    G2108_o2 <= 1'b0;
    G1126_o2 <= 1'b0;
    G1899_o2 <= 1'b0;
    G2134_o2 <= 1'b0;
    G1852_o2 <= 1'b0;
    G2116_o2 <= 1'b0;
    G2543_o2 <= 1'b0;
    G2727_o2 <= 1'b0;
    G2715_o2 <= 1'b0;
    G2832_o2 <= 1'b0;
    G1873_o2 <= 1'b0;
    G3291_o2 <= 1'b0;
    G5025_o2 <= 1'b0;
    G5036_o2 <= 1'b0;
    G3132_o2 <= 1'b0;
    G5038_o2 <= 1'b0;
    G5039_o2 <= 1'b0;
    n3118_inv <= 1'b0;
    n3121_inv <= 1'b0;
    n3124_inv <= 1'b0;
    n3127_inv <= 1'b0;
    n3984_lo_buf_o2 <= 1'b0;
    G1802_o2 <= 1'b0;
    G1804_o2 <= 1'b0;
    G1849_o2 <= 1'b0;
    G1851_o2 <= 1'b0;
    G2492_o2 <= 1'b0;
    G1799_o2 <= 1'b0;
    G4231_o2 <= 1'b0;
    G4234_o2 <= 1'b0;
    G4245_o2 <= 1'b0;
    G4247_o2 <= 1'b0;
    G1894_o2 <= 1'b0;
    G1846_o2 <= 1'b0;
    G4238_o2 <= 1'b0;
    G4249_o2 <= 1'b0;
    G2293_o2 <= 1'b0;
    G5022_o2 <= 1'b0;
    G5006_o2 <= 1'b0;
    G4944_o2 <= 1'b0;
    G4946_o2 <= 1'b0;
    G4954_o2 <= 1'b0;
    G4956_o2 <= 1'b0;
    G3546_o2 <= 1'b0;
    G3658_o2 <= 1'b0;
    G1344_o2 <= 1'b0;
    G2921_o2 <= 1'b0;
    n3912_lo_buf_o2 <= 1'b0;
    G1835_o2 <= 1'b0;
    G3810_o2 <= 1'b0;
    G3866_o2 <= 1'b0;
    G3811_o2 <= 1'b0;
    G2269_o2 <= 1'b0;
    G3812_o2 <= 1'b0;
    G3867_o2 <= 1'b0;
    G3868_o2 <= 1'b0;
    G3809_o2 <= 1'b0;
    G3716_o2 <= 1'b0;
    G4529_o2 <= 1'b0;
    G4670_o2 <= 1'b0;
    G4493_o2 <= 1'b0;
    G4580_o2 <= 1'b0;
    G3822_o2 <= 1'b0;
    G3877_o2 <= 1'b0;
    G4131_o2 <= 1'b0;
    G4170_o2 <= 1'b0;
    G4051_o2 <= 1'b0;
    G4065_o2 <= 1'b0;
    G4697_o2 <= 1'b0;
    G4706_o2 <= 1'b0;
    G2460_o2 <= 1'b0;
    G2454_o2 <= 1'b0;
    G2392_o2 <= 1'b0;
    G2386_o2 <= 1'b0;
    n4260_lo_buf_o2 <= 1'b0;
    n4272_lo_buf_o2 <= 1'b0;
    n4392_lo_buf_o2 <= 1'b0;
    n4404_lo_buf_o2 <= 1'b0;
    G1512_o2 <= 1'b0;
    G3135_o2 <= 1'b0;
    G2379_o2 <= 1'b0;
    n4164_lo_buf_o2 <= 1'b0;
    n4176_lo_buf_o2 <= 1'b0;
    n4224_lo_buf_o2 <= 1'b0;
    G2975_o2 <= 1'b0;
    G2978_o2 <= 1'b0;
    G2933_o2 <= 1'b0;
    G2936_o2 <= 1'b0;
    G1356_o2 <= 1'b0;
    G1359_o2 <= 1'b0;
    G1398_o2 <= 1'b0;
    G1401_o2 <= 1'b0;
  end
endmodule


