// Benchmark "c432" written by ABC on Sun Oct 29 19:31:46 2023

module c432 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36,
    G426, G427, G428, G429, G430, G431, G432  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36;
  output G426, G427, G428, G429, G430, G431, G432;
  reg n205_lo, n208_lo, n211_lo, n214_lo, n217_lo, n220_lo, n223_lo,
    n226_lo, n229_lo, n232_lo, n235_lo, n238_lo, n241_lo, n244_lo, n247_lo,
    n250_lo, n253_lo, n256_lo, n259_lo, n262_lo, n265_lo, n268_lo, n271_lo,
    n274_lo, n277_lo, n280_lo, n283_lo, n286_lo, n289_lo, n292_lo, n295_lo,
    n298_lo, n301_lo, n304_lo, n307_lo, n310_lo, n313_lo, n316_lo, n319_lo,
    n322_lo, n325_lo, n328_lo, n331_lo, n334_lo, n337_lo, n340_lo, n343_lo,
    n346_lo, n349_lo, n352_lo, n355_lo, n358_lo, n361_lo, n364_lo, n367_lo,
    n370_lo, n373_lo, n376_lo, n379_lo, n382_lo, n385_lo, n388_lo, n391_lo,
    n394_lo, n397_lo, n400_lo, n403_lo, n406_lo, n409_lo, n412_lo, n415_lo,
    n418_lo, n421_lo, n424_lo, n427_lo, n430_lo, n433_lo, n436_lo, n439_lo,
    n442_lo, n445_lo, n448_lo, n451_lo, n454_lo, n457_lo, n460_lo, n463_lo,
    n466_lo, n469_lo, n472_lo, n475_lo, n478_lo, n481_lo, n484_lo, n487_lo,
    n490_lo, n493_lo, n496_lo, n499_lo, n502_lo, n505_lo, n508_lo, n511_lo,
    n514_lo, n517_lo, n520_lo, n523_lo, n526_lo, n529_lo, n532_lo, n535_lo,
    n538_lo, n541_lo, n544_lo, n547_lo, n550_lo, n553_lo, n556_lo, n559_lo,
    n562_lo, n565_lo, n568_lo, n571_lo, n574_lo, n577_lo, n580_lo, n583_lo,
    n586_lo, n589_lo, n592_lo, n595_lo, n598_lo, n601_lo, n604_lo, n607_lo,
    n610_lo, n613_lo, n616_lo, n619_lo, n622_lo, n625_lo, n628_lo, n631_lo,
    n634_lo;
  wire new_G118_, new_G119_, new_G122_, new_G123_, new_G126_, new_G127_,
    new_G130_, new_G131_, new_G134_, new_G135_, new_G138_, new_G139_,
    new_G142_, new_G143_, new_G146_, new_G147_, new_G150_, new_G151_,
    new_G154_, new_G157_, new_G158_, new_G159_, new_G162_, new_G165_,
    new_G168_, new_G171_, new_G174_, new_G177_, new_G180_, new_G183_,
    new_G184_, new_G185_, new_G186_, new_G187_, new_G188_, new_G189_,
    new_G190_, new_G191_, new_G192_, new_G193_, new_G194_, new_G195_,
    new_G196_, new_G197_, new_G198_, new_G199_, new_G203_, new_G213_,
    new_G223_, new_G226_, new_G229_, new_G232_, new_G235_, new_G238_,
    new_G241_, new_G242_, new_G245_, new_G246_, new_G249_, new_G250_,
    new_G253_, new_G254_, new_G255_, new_G256_, new_G257_, new_G258_,
    new_G259_, new_G262_, new_G263_, new_G266_, new_G269_, new_G272_,
    new_G275_, new_G278_, new_G281_, new_G284_, new_G287_, new_G288_,
    new_G289_, new_G290_, new_G291_, new_G292_, new_G293_, new_G294_,
    new_G295_, new_G299_, new_G300_, new_G301_, new_G302_, new_G303_,
    new_G304_, new_G305_, new_G306_, new_G307_, new_G308_, new_G318_,
    new_G328_, new_G329_, new_G330_, new_G331_, new_G332_, new_G333_,
    new_G334_, new_G335_, new_G336_, new_G337_, new_G338_, new_G339_,
    new_G340_, new_G341_, new_G342_, new_G343_, new_G344_, new_G345_,
    new_G346_, new_G347_, new_G348_, new_G349_, new_G350_, new_G351_,
    new_G352_, new_G353_, new_G354_, new_G355_, new_G358_, new_G368_,
    new_G369_, new_G370_, new_G371_, new_G372_, new_G373_, new_G374_,
    new_G375_, new_G376_, new_G377_, new_G378_, new_G383_, new_G390_,
    new_G396_, new_G401_, new_G404_, new_G408_, new_G411_, new_G412_,
    new_G413_, new_G414_, new_G415_, new_G416_, new_G417_, new_G418_,
    new_G421_, new_G424_, new_G425_, n205_li, n208_li, n211_li, n214_li,
    n217_li, n220_li, n223_li, n226_li, n229_li, n232_li, n235_li, n238_li,
    n241_li, n244_li, n247_li, n250_li, n253_li, n256_li, n259_li, n262_li,
    n265_li, n268_li, n271_li, n274_li, n277_li, n280_li, n283_li, n286_li,
    n289_li, n292_li, n295_li, n298_li, n301_li, n304_li, n307_li, n310_li,
    n313_li, n316_li, n319_li, n322_li, n325_li, n328_li, n331_li, n334_li,
    n337_li, n340_li, n343_li, n346_li, n349_li, n352_li, n355_li, n358_li,
    n361_li, n364_li, n367_li, n370_li, n373_li, n376_li, n379_li, n382_li,
    n385_li, n388_li, n391_li, n394_li, n397_li, n400_li, n403_li, n406_li,
    n409_li, n412_li, n415_li, n418_li, n421_li, n424_li, n427_li, n430_li,
    n433_li, n436_li, n439_li, n442_li, n445_li, n448_li, n451_li, n454_li,
    n457_li, n460_li, n463_li, n466_li, n469_li, n472_li, n475_li, n478_li,
    n481_li, n484_li, n487_li, n490_li, n493_li, n496_li, n499_li, n502_li,
    n505_li, n508_li, n511_li, n514_li, n517_li, n520_li, n523_li, n526_li,
    n529_li, n532_li, n535_li, n538_li, n541_li, n544_li, n547_li, n550_li,
    n553_li, n556_li, n559_li, n562_li, n565_li, n568_li, n571_li, n574_li,
    n577_li, n580_li, n583_li, n586_li, n589_li, n592_li, n595_li, n598_li,
    n601_li, n604_li, n607_li, n610_li, n613_li, n616_li, n619_li, n622_li,
    n625_li, n628_li, n631_li, n634_li;
  assign new_G118_ = ~n214_lo;
  assign new_G119_ = ~n226_lo;
  assign new_G122_ = ~n250_lo;
  assign new_G123_ = ~n274_lo;
  assign new_G126_ = ~n298_lo;
  assign new_G127_ = ~n322_lo;
  assign new_G130_ = ~n346_lo;
  assign new_G131_ = ~n370_lo;
  assign new_G134_ = ~n394_lo;
  assign new_G135_ = ~n418_lo;
  assign new_G138_ = ~n442_lo;
  assign new_G139_ = ~n466_lo;
  assign new_G142_ = ~n490_lo;
  assign new_G143_ = ~n514_lo;
  assign new_G146_ = ~n538_lo;
  assign new_G147_ = ~n562_lo;
  assign new_G150_ = ~n586_lo;
  assign new_G151_ = ~n610_lo;
  assign new_G154_ = ~new_G118_ | ~n226_lo;
  assign new_G157_ = ~n238_lo & ~new_G119_;
  assign new_G158_ = ~n262_lo & ~new_G119_;
  assign new_G159_ = ~new_G122_ | ~n274_lo;
  assign new_G162_ = ~new_G126_ | ~n322_lo;
  assign new_G165_ = ~new_G130_ | ~n370_lo;
  assign new_G168_ = ~new_G134_ | ~n418_lo;
  assign new_G171_ = ~new_G138_ | ~n466_lo;
  assign new_G174_ = ~new_G142_ | ~n514_lo;
  assign new_G177_ = ~new_G146_ | ~n562_lo;
  assign new_G180_ = ~new_G150_ | ~n610_lo;
  assign new_G183_ = ~n286_lo & ~new_G123_;
  assign new_G184_ = ~n310_lo & ~new_G123_;
  assign new_G185_ = ~n334_lo & ~new_G127_;
  assign new_G186_ = ~n358_lo & ~new_G127_;
  assign new_G187_ = ~n382_lo & ~new_G131_;
  assign new_G188_ = ~n406_lo & ~new_G131_;
  assign new_G189_ = ~n430_lo & ~new_G135_;
  assign new_G190_ = ~n454_lo & ~new_G135_;
  assign new_G191_ = ~n478_lo & ~new_G139_;
  assign new_G192_ = ~n502_lo & ~new_G139_;
  assign new_G193_ = ~n526_lo & ~new_G143_;
  assign new_G194_ = ~n550_lo & ~new_G143_;
  assign new_G195_ = ~n574_lo & ~new_G147_;
  assign new_G196_ = ~n598_lo & ~new_G147_;
  assign new_G197_ = ~n622_lo & ~new_G151_;
  assign new_G198_ = ~n634_lo & ~new_G151_;
  assign new_G199_ = new_G180_ & new_G177_ & new_G174_ & new_G171_ & new_G168_ & new_G165_ & new_G154_ & new_G159_ & new_G162_;
  assign new_G203_ = ~new_G199_;
  assign new_G213_ = ~new_G199_;
  assign new_G223_ = new_G203_ ^ new_G154_;
  assign new_G226_ = new_G203_ ^ new_G159_;
  assign new_G229_ = new_G203_ ^ new_G162_;
  assign new_G232_ = new_G203_ ^ new_G165_;
  assign new_G235_ = new_G203_ ^ new_G168_;
  assign new_G238_ = new_G203_ ^ new_G171_;
  assign new_G241_ = ~n214_lo | ~new_G213_;
  assign new_G242_ = new_G203_ ^ new_G174_;
  assign new_G245_ = ~new_G213_ | ~n250_lo;
  assign new_G246_ = new_G203_ ^ new_G177_;
  assign new_G249_ = ~new_G213_ | ~n298_lo;
  assign new_G250_ = new_G203_ ^ new_G180_;
  assign new_G253_ = ~new_G213_ | ~n346_lo;
  assign new_G254_ = ~new_G213_ | ~n394_lo;
  assign new_G255_ = ~new_G213_ | ~n442_lo;
  assign new_G256_ = ~new_G213_ | ~n490_lo;
  assign new_G257_ = ~new_G213_ | ~n538_lo;
  assign new_G258_ = ~new_G213_ | ~n586_lo;
  assign new_G259_ = ~new_G223_ | ~new_G157_;
  assign new_G262_ = ~new_G223_ | ~new_G158_;
  assign new_G263_ = ~new_G226_ | ~new_G183_;
  assign new_G266_ = ~new_G229_ | ~new_G185_;
  assign new_G269_ = ~new_G232_ | ~new_G187_;
  assign new_G272_ = ~new_G235_ | ~new_G189_;
  assign new_G275_ = ~new_G238_ | ~new_G191_;
  assign new_G278_ = ~new_G242_ | ~new_G193_;
  assign new_G281_ = ~new_G246_ | ~new_G195_;
  assign new_G284_ = ~new_G250_ | ~new_G197_;
  assign new_G287_ = ~new_G226_ | ~new_G184_;
  assign new_G288_ = ~new_G229_ | ~new_G186_;
  assign new_G289_ = ~new_G232_ | ~new_G188_;
  assign new_G290_ = ~new_G235_ | ~new_G190_;
  assign new_G291_ = ~new_G238_ | ~new_G192_;
  assign new_G292_ = ~new_G242_ | ~new_G194_;
  assign new_G293_ = ~new_G246_ | ~new_G196_;
  assign new_G294_ = ~new_G250_ | ~new_G198_;
  assign new_G295_ = new_G284_ & new_G281_ & new_G278_ & new_G275_ & new_G272_ & new_G269_ & new_G259_ & new_G263_ & new_G266_;
  assign new_G299_ = ~new_G262_;
  assign new_G300_ = ~new_G287_;
  assign new_G301_ = ~new_G288_;
  assign new_G302_ = ~new_G289_;
  assign new_G303_ = ~new_G290_;
  assign new_G304_ = ~new_G291_;
  assign new_G305_ = ~new_G292_;
  assign new_G306_ = ~new_G293_;
  assign new_G307_ = ~new_G294_;
  assign new_G308_ = ~new_G295_;
  assign new_G318_ = ~new_G295_;
  assign new_G328_ = new_G308_ ^ new_G259_;
  assign new_G329_ = new_G308_ ^ new_G263_;
  assign new_G330_ = new_G308_ ^ new_G266_;
  assign new_G331_ = new_G308_ ^ new_G269_;
  assign new_G332_ = ~n238_lo | ~new_G318_;
  assign new_G333_ = new_G308_ ^ new_G272_;
  assign new_G334_ = ~new_G318_ | ~n286_lo;
  assign new_G335_ = new_G308_ ^ new_G275_;
  assign new_G336_ = ~new_G318_ | ~n334_lo;
  assign new_G337_ = new_G308_ ^ new_G278_;
  assign new_G338_ = ~new_G318_ | ~n382_lo;
  assign new_G339_ = new_G308_ ^ new_G281_;
  assign new_G340_ = ~new_G318_ | ~n430_lo;
  assign new_G341_ = new_G308_ ^ new_G284_;
  assign new_G342_ = ~new_G318_ | ~n478_lo;
  assign new_G343_ = ~new_G318_ | ~n526_lo;
  assign new_G344_ = ~new_G318_ | ~n574_lo;
  assign new_G345_ = ~new_G318_ | ~n622_lo;
  assign new_G346_ = ~new_G328_ | ~new_G299_;
  assign new_G347_ = ~new_G329_ | ~new_G300_;
  assign new_G348_ = ~new_G330_ | ~new_G301_;
  assign new_G349_ = ~new_G331_ | ~new_G302_;
  assign new_G350_ = ~new_G333_ | ~new_G303_;
  assign new_G351_ = ~new_G335_ | ~new_G304_;
  assign new_G352_ = ~new_G337_ | ~new_G305_;
  assign new_G353_ = ~new_G339_ | ~new_G306_;
  assign new_G354_ = ~new_G341_ | ~new_G307_;
  assign new_G355_ = new_G354_ & new_G353_ & new_G352_ & new_G351_ & new_G350_ & new_G349_ & new_G346_ & new_G347_ & new_G348_;
  assign new_G358_ = ~new_G355_;
  assign new_G368_ = ~n262_lo | ~new_G358_;
  assign new_G369_ = ~new_G358_ | ~n310_lo;
  assign new_G370_ = ~new_G358_ | ~n358_lo;
  assign new_G371_ = ~new_G358_ | ~n406_lo;
  assign new_G372_ = ~new_G358_ | ~n454_lo;
  assign new_G373_ = ~new_G358_ | ~n502_lo;
  assign new_G374_ = ~new_G358_ | ~n550_lo;
  assign new_G375_ = ~new_G358_ | ~n598_lo;
  assign new_G376_ = ~new_G358_ | ~n634_lo;
  assign new_G377_ = ~new_G368_ | ~n226_lo | ~new_G241_ | ~new_G332_;
  assign new_G378_ = ~n274_lo | ~new_G245_ | ~new_G334_ | ~new_G369_;
  assign new_G383_ = ~n322_lo | ~new_G249_ | ~new_G336_ | ~new_G370_;
  assign new_G390_ = ~n370_lo | ~new_G253_ | ~new_G338_ | ~new_G371_;
  assign new_G396_ = ~n418_lo | ~new_G254_ | ~new_G340_ | ~new_G372_;
  assign new_G401_ = ~n466_lo | ~new_G255_ | ~new_G342_ | ~new_G373_;
  assign new_G404_ = ~n514_lo | ~new_G256_ | ~new_G343_ | ~new_G374_;
  assign new_G408_ = ~n562_lo | ~new_G257_ | ~new_G344_ | ~new_G375_;
  assign new_G411_ = ~n610_lo | ~new_G258_ | ~new_G345_ | ~new_G376_;
  assign new_G412_ = ~new_G377_;
  assign new_G413_ = new_G411_ & new_G408_ & new_G404_ & new_G401_ & new_G396_ & new_G378_ & new_G383_ & new_G390_;
  assign new_G414_ = ~new_G390_;
  assign new_G415_ = ~new_G401_;
  assign new_G416_ = ~new_G404_;
  assign new_G417_ = ~new_G408_;
  assign new_G418_ = ~new_G383_ | ~new_G414_;
  assign new_G421_ = ~new_G396_ | ~new_G383_ | ~new_G390_ | ~new_G415_;
  assign new_G424_ = ~new_G396_ | ~new_G390_ | ~new_G416_;
  assign new_G425_ = ~new_G417_ | ~new_G383_ | ~new_G390_ | ~new_G404_;
  assign G426 = ~new_G199_;
  assign G427 = ~new_G295_;
  assign G428 = ~new_G355_;
  assign G429 = ~new_G412_ & ~new_G413_;
  assign G430 = ~new_G396_ | ~new_G378_ | ~new_G383_ | ~new_G418_;
  assign G431 = ~new_G424_ | ~new_G378_ | ~new_G383_ | ~new_G421_;
  assign G432 = ~new_G425_ | ~new_G378_ | ~new_G418_ | ~new_G421_;
  assign n205_li = G1;
  assign n208_li = n205_lo;
  assign n211_li = n208_lo;
  assign n214_li = n211_lo;
  assign n217_li = G2;
  assign n220_li = n217_lo;
  assign n223_li = n220_lo;
  assign n226_li = n223_lo;
  assign n229_li = G3;
  assign n232_li = n229_lo;
  assign n235_li = n232_lo;
  assign n238_li = n235_lo;
  assign n241_li = G4;
  assign n244_li = n241_lo;
  assign n247_li = n244_lo;
  assign n250_li = n247_lo;
  assign n253_li = G5;
  assign n256_li = n253_lo;
  assign n259_li = n256_lo;
  assign n262_li = n259_lo;
  assign n265_li = G6;
  assign n268_li = n265_lo;
  assign n271_li = n268_lo;
  assign n274_li = n271_lo;
  assign n277_li = G7;
  assign n280_li = n277_lo;
  assign n283_li = n280_lo;
  assign n286_li = n283_lo;
  assign n289_li = G8;
  assign n292_li = n289_lo;
  assign n295_li = n292_lo;
  assign n298_li = n295_lo;
  assign n301_li = G9;
  assign n304_li = n301_lo;
  assign n307_li = n304_lo;
  assign n310_li = n307_lo;
  assign n313_li = G10;
  assign n316_li = n313_lo;
  assign n319_li = n316_lo;
  assign n322_li = n319_lo;
  assign n325_li = G11;
  assign n328_li = n325_lo;
  assign n331_li = n328_lo;
  assign n334_li = n331_lo;
  assign n337_li = G12;
  assign n340_li = n337_lo;
  assign n343_li = n340_lo;
  assign n346_li = n343_lo;
  assign n349_li = G13;
  assign n352_li = n349_lo;
  assign n355_li = n352_lo;
  assign n358_li = n355_lo;
  assign n361_li = G14;
  assign n364_li = n361_lo;
  assign n367_li = n364_lo;
  assign n370_li = n367_lo;
  assign n373_li = G15;
  assign n376_li = n373_lo;
  assign n379_li = n376_lo;
  assign n382_li = n379_lo;
  assign n385_li = G16;
  assign n388_li = n385_lo;
  assign n391_li = n388_lo;
  assign n394_li = n391_lo;
  assign n397_li = G17;
  assign n400_li = n397_lo;
  assign n403_li = n400_lo;
  assign n406_li = n403_lo;
  assign n409_li = G18;
  assign n412_li = n409_lo;
  assign n415_li = n412_lo;
  assign n418_li = n415_lo;
  assign n421_li = G19;
  assign n424_li = n421_lo;
  assign n427_li = n424_lo;
  assign n430_li = n427_lo;
  assign n433_li = G20;
  assign n436_li = n433_lo;
  assign n439_li = n436_lo;
  assign n442_li = n439_lo;
  assign n445_li = G21;
  assign n448_li = n445_lo;
  assign n451_li = n448_lo;
  assign n454_li = n451_lo;
  assign n457_li = G22;
  assign n460_li = n457_lo;
  assign n463_li = n460_lo;
  assign n466_li = n463_lo;
  assign n469_li = G23;
  assign n472_li = n469_lo;
  assign n475_li = n472_lo;
  assign n478_li = n475_lo;
  assign n481_li = G24;
  assign n484_li = n481_lo;
  assign n487_li = n484_lo;
  assign n490_li = n487_lo;
  assign n493_li = G25;
  assign n496_li = n493_lo;
  assign n499_li = n496_lo;
  assign n502_li = n499_lo;
  assign n505_li = G26;
  assign n508_li = n505_lo;
  assign n511_li = n508_lo;
  assign n514_li = n511_lo;
  assign n517_li = G27;
  assign n520_li = n517_lo;
  assign n523_li = n520_lo;
  assign n526_li = n523_lo;
  assign n529_li = G28;
  assign n532_li = n529_lo;
  assign n535_li = n532_lo;
  assign n538_li = n535_lo;
  assign n541_li = G29;
  assign n544_li = n541_lo;
  assign n547_li = n544_lo;
  assign n550_li = n547_lo;
  assign n553_li = G30;
  assign n556_li = n553_lo;
  assign n559_li = n556_lo;
  assign n562_li = n559_lo;
  assign n565_li = G31;
  assign n568_li = n565_lo;
  assign n571_li = n568_lo;
  assign n574_li = n571_lo;
  assign n577_li = G32;
  assign n580_li = n577_lo;
  assign n583_li = n580_lo;
  assign n586_li = n583_lo;
  assign n589_li = G33;
  assign n592_li = n589_lo;
  assign n595_li = n592_lo;
  assign n598_li = n595_lo;
  assign n601_li = G34;
  assign n604_li = n601_lo;
  assign n607_li = n604_lo;
  assign n610_li = n607_lo;
  assign n613_li = G35;
  assign n616_li = n613_lo;
  assign n619_li = n616_lo;
  assign n622_li = n619_lo;
  assign n625_li = G36;
  assign n628_li = n625_lo;
  assign n631_li = n628_lo;
  assign n634_li = n631_lo;
  always @ (posedge clock) begin
    n205_lo <= n205_li;
    n208_lo <= n208_li;
    n211_lo <= n211_li;
    n214_lo <= n214_li;
    n217_lo <= n217_li;
    n220_lo <= n220_li;
    n223_lo <= n223_li;
    n226_lo <= n226_li;
    n229_lo <= n229_li;
    n232_lo <= n232_li;
    n235_lo <= n235_li;
    n238_lo <= n238_li;
    n241_lo <= n241_li;
    n244_lo <= n244_li;
    n247_lo <= n247_li;
    n250_lo <= n250_li;
    n253_lo <= n253_li;
    n256_lo <= n256_li;
    n259_lo <= n259_li;
    n262_lo <= n262_li;
    n265_lo <= n265_li;
    n268_lo <= n268_li;
    n271_lo <= n271_li;
    n274_lo <= n274_li;
    n277_lo <= n277_li;
    n280_lo <= n280_li;
    n283_lo <= n283_li;
    n286_lo <= n286_li;
    n289_lo <= n289_li;
    n292_lo <= n292_li;
    n295_lo <= n295_li;
    n298_lo <= n298_li;
    n301_lo <= n301_li;
    n304_lo <= n304_li;
    n307_lo <= n307_li;
    n310_lo <= n310_li;
    n313_lo <= n313_li;
    n316_lo <= n316_li;
    n319_lo <= n319_li;
    n322_lo <= n322_li;
    n325_lo <= n325_li;
    n328_lo <= n328_li;
    n331_lo <= n331_li;
    n334_lo <= n334_li;
    n337_lo <= n337_li;
    n340_lo <= n340_li;
    n343_lo <= n343_li;
    n346_lo <= n346_li;
    n349_lo <= n349_li;
    n352_lo <= n352_li;
    n355_lo <= n355_li;
    n358_lo <= n358_li;
    n361_lo <= n361_li;
    n364_lo <= n364_li;
    n367_lo <= n367_li;
    n370_lo <= n370_li;
    n373_lo <= n373_li;
    n376_lo <= n376_li;
    n379_lo <= n379_li;
    n382_lo <= n382_li;
    n385_lo <= n385_li;
    n388_lo <= n388_li;
    n391_lo <= n391_li;
    n394_lo <= n394_li;
    n397_lo <= n397_li;
    n400_lo <= n400_li;
    n403_lo <= n403_li;
    n406_lo <= n406_li;
    n409_lo <= n409_li;
    n412_lo <= n412_li;
    n415_lo <= n415_li;
    n418_lo <= n418_li;
    n421_lo <= n421_li;
    n424_lo <= n424_li;
    n427_lo <= n427_li;
    n430_lo <= n430_li;
    n433_lo <= n433_li;
    n436_lo <= n436_li;
    n439_lo <= n439_li;
    n442_lo <= n442_li;
    n445_lo <= n445_li;
    n448_lo <= n448_li;
    n451_lo <= n451_li;
    n454_lo <= n454_li;
    n457_lo <= n457_li;
    n460_lo <= n460_li;
    n463_lo <= n463_li;
    n466_lo <= n466_li;
    n469_lo <= n469_li;
    n472_lo <= n472_li;
    n475_lo <= n475_li;
    n478_lo <= n478_li;
    n481_lo <= n481_li;
    n484_lo <= n484_li;
    n487_lo <= n487_li;
    n490_lo <= n490_li;
    n493_lo <= n493_li;
    n496_lo <= n496_li;
    n499_lo <= n499_li;
    n502_lo <= n502_li;
    n505_lo <= n505_li;
    n508_lo <= n508_li;
    n511_lo <= n511_li;
    n514_lo <= n514_li;
    n517_lo <= n517_li;
    n520_lo <= n520_li;
    n523_lo <= n523_li;
    n526_lo <= n526_li;
    n529_lo <= n529_li;
    n532_lo <= n532_li;
    n535_lo <= n535_li;
    n538_lo <= n538_li;
    n541_lo <= n541_li;
    n544_lo <= n544_li;
    n547_lo <= n547_li;
    n550_lo <= n550_li;
    n553_lo <= n553_li;
    n556_lo <= n556_li;
    n559_lo <= n559_li;
    n562_lo <= n562_li;
    n565_lo <= n565_li;
    n568_lo <= n568_li;
    n571_lo <= n571_li;
    n574_lo <= n574_li;
    n577_lo <= n577_li;
    n580_lo <= n580_li;
    n583_lo <= n583_li;
    n586_lo <= n586_li;
    n589_lo <= n589_li;
    n592_lo <= n592_li;
    n595_lo <= n595_li;
    n598_lo <= n598_li;
    n601_lo <= n601_li;
    n604_lo <= n604_li;
    n607_lo <= n607_li;
    n610_lo <= n610_li;
    n613_lo <= n613_li;
    n616_lo <= n616_li;
    n619_lo <= n619_li;
    n622_lo <= n622_li;
    n625_lo <= n625_li;
    n628_lo <= n628_li;
    n631_lo <= n631_li;
    n634_lo <= n634_li;
  end
  initial begin
    n205_lo <= 1'b0;
    n208_lo <= 1'b0;
    n211_lo <= 1'b0;
    n214_lo <= 1'b0;
    n217_lo <= 1'b0;
    n220_lo <= 1'b0;
    n223_lo <= 1'b0;
    n226_lo <= 1'b0;
    n229_lo <= 1'b0;
    n232_lo <= 1'b0;
    n235_lo <= 1'b0;
    n238_lo <= 1'b0;
    n241_lo <= 1'b0;
    n244_lo <= 1'b0;
    n247_lo <= 1'b0;
    n250_lo <= 1'b0;
    n253_lo <= 1'b0;
    n256_lo <= 1'b0;
    n259_lo <= 1'b0;
    n262_lo <= 1'b0;
    n265_lo <= 1'b0;
    n268_lo <= 1'b0;
    n271_lo <= 1'b0;
    n274_lo <= 1'b0;
    n277_lo <= 1'b0;
    n280_lo <= 1'b0;
    n283_lo <= 1'b0;
    n286_lo <= 1'b0;
    n289_lo <= 1'b0;
    n292_lo <= 1'b0;
    n295_lo <= 1'b0;
    n298_lo <= 1'b0;
    n301_lo <= 1'b0;
    n304_lo <= 1'b0;
    n307_lo <= 1'b0;
    n310_lo <= 1'b0;
    n313_lo <= 1'b0;
    n316_lo <= 1'b0;
    n319_lo <= 1'b0;
    n322_lo <= 1'b0;
    n325_lo <= 1'b0;
    n328_lo <= 1'b0;
    n331_lo <= 1'b0;
    n334_lo <= 1'b0;
    n337_lo <= 1'b0;
    n340_lo <= 1'b0;
    n343_lo <= 1'b0;
    n346_lo <= 1'b0;
    n349_lo <= 1'b0;
    n352_lo <= 1'b0;
    n355_lo <= 1'b0;
    n358_lo <= 1'b0;
    n361_lo <= 1'b0;
    n364_lo <= 1'b0;
    n367_lo <= 1'b0;
    n370_lo <= 1'b0;
    n373_lo <= 1'b0;
    n376_lo <= 1'b0;
    n379_lo <= 1'b0;
    n382_lo <= 1'b0;
    n385_lo <= 1'b0;
    n388_lo <= 1'b0;
    n391_lo <= 1'b0;
    n394_lo <= 1'b0;
    n397_lo <= 1'b0;
    n400_lo <= 1'b0;
    n403_lo <= 1'b0;
    n406_lo <= 1'b0;
    n409_lo <= 1'b0;
    n412_lo <= 1'b0;
    n415_lo <= 1'b0;
    n418_lo <= 1'b0;
    n421_lo <= 1'b0;
    n424_lo <= 1'b0;
    n427_lo <= 1'b0;
    n430_lo <= 1'b0;
    n433_lo <= 1'b0;
    n436_lo <= 1'b0;
    n439_lo <= 1'b0;
    n442_lo <= 1'b0;
    n445_lo <= 1'b0;
    n448_lo <= 1'b0;
    n451_lo <= 1'b0;
    n454_lo <= 1'b0;
    n457_lo <= 1'b0;
    n460_lo <= 1'b0;
    n463_lo <= 1'b0;
    n466_lo <= 1'b0;
    n469_lo <= 1'b0;
    n472_lo <= 1'b0;
    n475_lo <= 1'b0;
    n478_lo <= 1'b0;
    n481_lo <= 1'b0;
    n484_lo <= 1'b0;
    n487_lo <= 1'b0;
    n490_lo <= 1'b0;
    n493_lo <= 1'b0;
    n496_lo <= 1'b0;
    n499_lo <= 1'b0;
    n502_lo <= 1'b0;
    n505_lo <= 1'b0;
    n508_lo <= 1'b0;
    n511_lo <= 1'b0;
    n514_lo <= 1'b0;
    n517_lo <= 1'b0;
    n520_lo <= 1'b0;
    n523_lo <= 1'b0;
    n526_lo <= 1'b0;
    n529_lo <= 1'b0;
    n532_lo <= 1'b0;
    n535_lo <= 1'b0;
    n538_lo <= 1'b0;
    n541_lo <= 1'b0;
    n544_lo <= 1'b0;
    n547_lo <= 1'b0;
    n550_lo <= 1'b0;
    n553_lo <= 1'b0;
    n556_lo <= 1'b0;
    n559_lo <= 1'b0;
    n562_lo <= 1'b0;
    n565_lo <= 1'b0;
    n568_lo <= 1'b0;
    n571_lo <= 1'b0;
    n574_lo <= 1'b0;
    n577_lo <= 1'b0;
    n580_lo <= 1'b0;
    n583_lo <= 1'b0;
    n586_lo <= 1'b0;
    n589_lo <= 1'b0;
    n592_lo <= 1'b0;
    n595_lo <= 1'b0;
    n598_lo <= 1'b0;
    n601_lo <= 1'b0;
    n604_lo <= 1'b0;
    n607_lo <= 1'b0;
    n610_lo <= 1'b0;
    n613_lo <= 1'b0;
    n616_lo <= 1'b0;
    n619_lo <= 1'b0;
    n622_lo <= 1'b0;
    n625_lo <= 1'b0;
    n628_lo <= 1'b0;
    n631_lo <= 1'b0;
    n634_lo <= 1'b0;
  end
endmodule


