// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:48 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479,
    G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491,
    G492, G493, G494, G495, G496, G497, G498, G499  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478,
    G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490,
    G491, G492, G493, G494, G495, G496, G497, G498, G499;
  reg n286_lo, n298_lo, n310_lo, n322_lo, n334_lo, n346_lo, n358_lo,
    n370_lo, n382_lo, n394_lo, n406_lo, n418_lo, n430_lo, n442_lo, n454_lo,
    n466_lo, n478_lo, n490_lo, n502_lo, n514_lo, n526_lo, n538_lo, n550_lo,
    n562_lo, n574_lo, n586_lo, n598_lo, n610_lo, n622_lo, n634_lo, n646_lo,
    n658_lo, n661_lo, n673_lo, n685_lo, n697_lo, n709_lo, n721_lo, n733_lo,
    n745_lo, n757_lo, n1248_o2, n1249_o2, n1250_o2, n1251_o2, n1252_o2,
    n1253_o2, n1254_o2, n1255_o2, n1207_o2, n1208_o2, n1209_o2, n1210_o2,
    n1211_o2, n1212_o2, n1213_o2, n1214_o2, n1215_o2, n1216_o2, n1217_o2,
    n1218_o2, n1219_o2, n1220_o2, n1221_o2, n1222_o2, n1223_o2, n1224_o2,
    n1225_o2, n1226_o2, n1227_o2, n1228_o2, n1229_o2, n1230_o2, n1231_o2,
    n1232_o2, n1233_o2, n1234_o2, n1235_o2, n1236_o2, n1237_o2, n1238_o2,
    G374_o2, G376_o2, G370_o2, G372_o2, G373_o2, G377_o2, G371_o2, G375_o2,
    G354_o2, G356_o2, G350_o2, G352_o2, G353_o2, G357_o2, G351_o2, G355_o2,
    G386_o2, G391_o2, n283_lo_buf_o2, n295_lo_buf_o2, n307_lo_buf_o2,
    n319_lo_buf_o2, n331_lo_buf_o2, n343_lo_buf_o2, n355_lo_buf_o2,
    n367_lo_buf_o2, n379_lo_buf_o2, n391_lo_buf_o2, n403_lo_buf_o2,
    n415_lo_buf_o2, n427_lo_buf_o2, n439_lo_buf_o2, n451_lo_buf_o2,
    n463_lo_buf_o2, n475_lo_buf_o2, n487_lo_buf_o2, n499_lo_buf_o2,
    n511_lo_buf_o2, n523_lo_buf_o2, n535_lo_buf_o2, n547_lo_buf_o2,
    n559_lo_buf_o2, n571_lo_buf_o2, n583_lo_buf_o2, n595_lo_buf_o2,
    n607_lo_buf_o2, n619_lo_buf_o2, n631_lo_buf_o2, n643_lo_buf_o2,
    n655_lo_buf_o2, G234_o2, G247_o2, G260_o2, G273_o2, G286_o2, G299_o2,
    G312_o2, G325_o2, n667_lo_buf_o2, n679_lo_buf_o2, n691_lo_buf_o2,
    n703_lo_buf_o2, n715_lo_buf_o2, n727_lo_buf_o2, n739_lo_buf_o2,
    n751_lo_buf_o2, n763_lo_buf_o2, G186_o2, G189_o2, G192_o2, G195_o2,
    G198_o2, G201_o2, G204_o2, G207_o2, n280_lo_buf_o2, n292_lo_buf_o2,
    n304_lo_buf_o2, n316_lo_buf_o2, n328_lo_buf_o2, n340_lo_buf_o2,
    n352_lo_buf_o2, n364_lo_buf_o2, n376_lo_buf_o2, n388_lo_buf_o2,
    n400_lo_buf_o2, n412_lo_buf_o2, n424_lo_buf_o2, n436_lo_buf_o2,
    n448_lo_buf_o2, n460_lo_buf_o2, n472_lo_buf_o2, n484_lo_buf_o2,
    n496_lo_buf_o2, n508_lo_buf_o2, n520_lo_buf_o2, n532_lo_buf_o2,
    n544_lo_buf_o2, n556_lo_buf_o2, n568_lo_buf_o2, n580_lo_buf_o2,
    n592_lo_buf_o2, n604_lo_buf_o2, n616_lo_buf_o2, n628_lo_buf_o2,
    n640_lo_buf_o2, n652_lo_buf_o2;
  wire new_new_n451__, new_new_n453__, new_new_n455__, new_new_n457__,
    new_new_n459__, new_new_n461__, new_new_n463__, new_new_n465__,
    new_new_n467__, new_new_n469__, new_new_n471__, new_new_n473__,
    new_new_n475__, new_new_n477__, new_new_n479__, new_new_n481__,
    new_new_n483__, new_new_n485__, new_new_n487__, new_new_n489__,
    new_new_n491__, new_new_n493__, new_new_n495__, new_new_n497__,
    new_new_n499__, new_new_n501__, new_new_n503__, new_new_n505__,
    new_new_n507__, new_new_n509__, new_new_n511__, new_new_n513__,
    new_new_n515__, new_new_n517__, new_new_n519__, new_new_n521__,
    new_new_n523__, new_new_n525__, new_new_n527__, new_new_n529__,
    new_new_n531__, new_new_n532__, new_new_n533__, new_new_n534__,
    new_new_n535__, new_new_n536__, new_new_n537__, new_new_n538__,
    new_new_n539__, new_new_n540__, new_new_n541__, new_new_n542__,
    new_new_n543__, new_new_n544__, new_new_n545__, new_new_n546__,
    new_new_n547__, new_new_n548__, new_new_n549__, new_new_n550__,
    new_new_n551__, new_new_n552__, new_new_n553__, new_new_n554__,
    new_new_n555__, new_new_n556__, new_new_n557__, new_new_n558__,
    new_new_n559__, new_new_n560__, new_new_n561__, new_new_n562__,
    new_new_n563__, new_new_n564__, new_new_n565__, new_new_n566__,
    new_new_n567__, new_new_n568__, new_new_n569__, new_new_n570__,
    new_new_n571__, new_new_n572__, new_new_n573__, new_new_n574__,
    new_new_n575__, new_new_n576__, new_new_n577__, new_new_n578__,
    new_new_n579__, new_new_n580__, new_new_n581__, new_new_n582__,
    new_new_n583__, new_new_n584__, new_new_n585__, new_new_n586__,
    new_new_n587__, new_new_n588__, new_new_n589__, new_new_n590__,
    new_new_n591__, new_new_n592__, new_new_n593__, new_new_n594__,
    new_new_n595__, new_new_n597__, new_new_n599__, new_new_n601__,
    new_new_n603__, new_new_n605__, new_new_n607__, new_new_n609__,
    new_new_n611__, new_new_n613__, new_new_n614__, new_new_n615__,
    new_new_n616__, new_new_n617__, new_new_n618__, new_new_n619__,
    new_new_n620__, new_new_n621__, new_new_n622__, new_new_n623__,
    new_new_n624__, new_new_n625__, new_new_n626__, new_new_n627__,
    new_new_n628__, new_new_n629__, new_new_n631__, new_new_n633__,
    new_new_n635__, new_new_n637__, new_new_n639__, new_new_n641__,
    new_new_n643__, new_new_n645__, new_new_n647__, new_new_n649__,
    new_new_n651__, new_new_n653__, new_new_n655__, new_new_n657__,
    new_new_n659__, new_new_n661__, new_new_n663__, new_new_n665__,
    new_new_n667__, new_new_n669__, new_new_n671__, new_new_n673__,
    new_new_n675__, new_new_n677__, new_new_n679__, new_new_n681__,
    new_new_n683__, new_new_n685__, new_new_n687__, new_new_n689__,
    new_new_n691__, new_new_n693__, new_new_n694__, new_new_n695__,
    new_new_n696__, new_new_n697__, new_new_n698__, new_new_n699__,
    new_new_n700__, new_new_n701__, new_new_n702__, new_new_n703__,
    new_new_n704__, new_new_n705__, new_new_n706__, new_new_n707__,
    new_new_n708__, new_new_n709__, new_new_n710__, new_new_n711__,
    new_new_n712__, new_new_n713__, new_new_n714__, new_new_n715__,
    new_new_n716__, new_new_n717__, new_new_n718__, new_new_n719__,
    new_new_n720__, new_new_n721__, new_new_n722__, new_new_n723__,
    new_new_n724__, new_new_n725__, new_new_n726__, new_new_n727__,
    new_new_n728__, new_new_n729__, new_new_n730__, new_new_n731__,
    new_new_n732__, new_new_n733__, new_new_n734__, new_new_n735__,
    new_new_n736__, new_new_n737__, new_new_n738__, new_new_n739__,
    new_new_n740__, new_new_n741__, new_new_n742__, new_new_n743__,
    new_new_n744__, new_new_n745__, new_new_n746__, new_new_n747__,
    new_new_n748__, new_new_n749__, new_new_n750__, new_new_n751__,
    new_new_n752__, new_new_n753__, new_new_n754__, new_new_n755__,
    new_new_n756__, new_new_n757__, new_new_n758__, new_new_n759__,
    new_new_n760__, new_new_n761__, new_new_n762__, new_new_n763__,
    new_new_n764__, new_new_n765__, new_new_n766__, new_new_n767__,
    new_new_n768__, new_new_n769__, new_new_n770__, new_new_n771__,
    new_new_n772__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n786__, new_new_n787__,
    new_new_n788__, new_new_n789__, new_new_n790__, new_new_n791__,
    new_new_n792__, new_new_n793__, new_new_n794__, new_new_n795__,
    new_new_n796__, new_new_n797__, new_new_n798__, new_new_n799__,
    new_new_n800__, new_new_n801__, new_new_n802__, new_new_n803__,
    new_new_n804__, new_new_n805__, new_new_n806__, new_new_n807__,
    new_new_n808__, new_new_n809__, new_new_n810__, new_new_n811__,
    new_new_n812__, new_new_n813__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n850__, new_new_n851__,
    new_new_n852__, new_new_n853__, new_new_n854__, new_new_n855__,
    new_new_n856__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n864__, new_new_n865__, new_new_n866__, new_new_n867__,
    new_new_n868__, new_new_n869__, new_new_n870__, new_new_n871__,
    new_new_n872__, new_new_n873__, new_new_n874__, new_new_n875__,
    new_new_n876__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n880__, new_new_n881__, new_new_n882__, new_new_n883__,
    new_new_n884__, new_new_n885__, new_new_n886__, new_new_n887__,
    new_new_n888__, new_new_n889__, new_new_n890__, new_new_n891__,
    new_new_n892__, new_new_n893__, new_new_n894__, new_new_n895__,
    new_new_n896__, new_new_n897__, new_new_n898__, new_new_n899__,
    new_new_n900__, new_new_n901__, new_new_n902__, new_new_n903__,
    new_new_n904__, new_new_n905__, new_new_n906__, new_new_n907__,
    new_new_n908__, new_new_n909__, new_new_n910__, new_new_n911__,
    new_new_n912__, new_new_n913__, new_new_n914__, new_new_n915__,
    new_new_n916__, new_new_n917__, new_new_n918__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n966__, new_new_n967__,
    new_new_n968__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n987__,
    new_new_n988__, new_new_n989__, new_new_n990__, new_new_n991__,
    new_new_n992__, new_new_n993__, new_new_n994__, new_new_n995__,
    new_new_n996__, new_new_n997__, new_new_n998__, new_new_n999__,
    new_new_n1000__, new_new_n1001__, new_new_n1002__, new_new_n1003__,
    new_new_n1004__, new_new_n1005__, new_new_n1006__, new_new_n1007__,
    new_new_n1008__, new_new_n1009__, new_new_n1010__, new_new_n1011__,
    new_new_n1012__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1022__, new_new_n1023__,
    new_new_n1024__, new_new_n1025__, new_new_n1026__, new_new_n1027__,
    new_new_n1028__, new_new_n1029__, new_new_n1030__, new_new_n1031__,
    new_new_n1032__, new_new_n1033__, new_new_n1034__, new_new_n1035__,
    new_new_n1036__, new_new_n1037__, new_new_n1038__, new_new_n1039__,
    new_new_n1040__, new_new_n1041__, new_new_n1042__, new_new_n1043__,
    new_new_n1044__, new_new_n1045__, new_new_n1046__, new_new_n1047__,
    new_new_n1048__, new_new_n1049__, new_new_n1050__, new_new_n1051__,
    new_new_n1052__, new_new_n1053__, new_new_n1054__, new_new_n1055__,
    new_new_n1056__, new_new_n1057__, new_new_n1058__, new_new_n1059__,
    new_new_n1060__, new_new_n1061__, new_new_n1062__, new_new_n1063__,
    new_new_n1064__, new_new_n1065__, new_new_n1066__, new_new_n1067__,
    new_new_n1068__, new_new_n1069__, new_new_n1070__, new_new_n1071__,
    new_new_n1072__, new_new_n1073__, new_new_n1074__, new_new_n1075__,
    new_new_n1076__, new_new_n1077__, new_new_n1078__, new_new_n1079__,
    new_new_n1080__, new_new_n1081__, new_new_n1082__, new_new_n1083__,
    new_new_n1084__, new_new_n1085__, new_new_n1086__, new_new_n1087__,
    new_new_n1088__, new_new_n1089__, new_new_n1090__, new_new_n1091__,
    new_new_n1092__, new_new_n1093__, new_new_n1094__, new_new_n1095__,
    new_new_n1096__, new_new_n1097__, new_new_n1098__, new_new_n1099__,
    new_new_n1100__, new_new_n1101__, new_new_n1102__, new_new_n1103__,
    new_new_n1104__, new_new_n1105__, new_new_n1106__, new_new_n1107__,
    new_new_n1108__, new_new_n1109__, new_new_n1110__, new_new_n1111__,
    new_new_n1112__, new_new_n1113__, new_new_n1114__, new_new_n1115__,
    new_new_n1116__, new_new_n1117__, new_new_n1118__, new_new_n1119__,
    new_new_n1120__, new_new_n1121__, new_new_n1122__, new_new_n1123__,
    new_new_n1124__, new_new_n1125__, new_new_n1126__, new_new_n1127__,
    new_new_n1128__, new_new_n1129__, new_new_n1130__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1142__, new_new_n1143__,
    new_new_n1144__, new_new_n1145__, new_new_n1146__, new_new_n1147__,
    new_new_n1148__, new_new_n1149__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1170__, new_new_n1171__,
    new_new_n1172__, new_new_n1173__, new_new_n1174__, new_new_n1175__,
    new_new_n1176__, new_new_n1177__, new_new_n1178__, new_new_n1179__,
    new_new_n1180__, new_new_n1181__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1202__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1206__, new_new_n1207__,
    new_new_n1208__, new_new_n1209__, new_new_n1210__, new_new_n1211__,
    new_new_n1212__, new_new_n1213__, new_new_n1214__, new_new_n1215__,
    new_new_n1216__, new_new_n1217__, new_new_n1218__, new_new_n1219__,
    new_new_n1220__, new_new_n1221__, new_new_n1222__, new_new_n1223__,
    new_new_n1224__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1232__, new_new_n1233__, new_new_n1234__, new_new_n1235__,
    new_new_n1236__, new_new_n1237__, new_new_n1238__, new_new_n1239__,
    new_new_n1240__, new_new_n1241__, new_new_n1242__, new_new_n1243__,
    new_new_n1244__, new_new_n1245__, new_new_n1246__, new_new_n1247__,
    new_new_n1248__, new_new_n1249__, new_new_n1250__, new_new_n1251__,
    new_new_n1252__, new_new_n1253__, new_new_n1254__, new_new_n1255__,
    new_new_n1256__, new_new_n1257__, new_new_n1258__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1265__, new_new_n1266__, new_new_n1267__,
    new_new_n1268__, new_new_n1269__, new_new_n1270__, new_new_n1271__,
    new_new_n1272__, new_new_n1273__, new_new_n1274__, new_new_n1275__,
    new_new_n1276__, new_new_n1277__, new_new_n1278__, new_new_n1279__,
    new_new_n1280__, new_new_n1281__, new_new_n1282__, new_new_n1283__,
    new_new_n1284__, new_new_n1285__, new_new_n1286__, new_new_n1287__,
    new_new_n1288__, new_new_n1289__, new_new_n1290__, new_new_n1291__,
    new_new_n1292__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1319__,
    new_new_n1320__, new_new_n1321__, new_new_n1322__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1336__, new_new_n1337__, new_new_n1338__, new_new_n1339__,
    new_new_n1340__, new_new_n1341__, new_new_n1342__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1346__, new_new_n1347__,
    new_new_n1348__, new_new_n1349__, new_new_n1350__, new_new_n1351__,
    new_new_n1352__, new_new_n1353__, new_new_n1354__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1362__, new_new_n1363__,
    new_new_n1364__, new_new_n1365__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1369__, new_new_n1370__, new_new_n1371__,
    new_new_n1372__, new_new_n1373__, new_new_n1374__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1394__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1482__, new_new_n1483__,
    new_new_n1484__, new_new_n1485__, new_new_n1486__, new_new_n1487__,
    new_new_n1488__, new_new_n1489__, new_new_n1490__, new_new_n1491__,
    new_new_n1492__, new_new_n1493__, new_new_n1494__, new_new_n1495__,
    new_new_n1496__, new_new_n1497__, new_new_n1498__, new_new_n1499__,
    new_new_n1500__, new_new_n1501__, new_new_n1502__, new_new_n1503__,
    new_new_n1504__, new_new_n1505__, new_new_n1506__, new_new_n1507__,
    new_new_n1508__, new_new_n1509__, new_new_n1510__, new_new_n1511__,
    new_new_n1512__, new_new_n1513__, new_new_n1514__, new_new_n1515__,
    new_new_n1516__, new_new_n1517__, new_new_n1518__, new_new_n1519__,
    new_new_n1520__, new_new_n1521__, new_new_n1522__, new_new_n1523__,
    new_new_n1524__, new_new_n1525__, new_new_n1526__, new_new_n1527__,
    new_new_n1528__, new_new_n1529__, new_new_n1530__, new_new_n1531__,
    new_new_n1532__, new_new_n1533__, new_new_n1534__, new_new_n1535__,
    new_new_n1536__, new_new_n1537__, new_new_n1538__, new_new_n1539__,
    new_new_n1540__, new_new_n1541__, new_new_n1542__, new_new_n1543__,
    new_new_n1544__, new_new_n1545__, new_new_n1546__, new_new_n1547__,
    new_new_n1548__, new_new_n1549__, new_new_n1550__, new_new_n1551__,
    new_new_n1552__, new_new_n1553__, new_new_n1554__, new_new_n1555__,
    new_new_n1556__, new_new_n1557__, new_new_n1558__, new_new_n1559__,
    new_new_n1780__, new_new_n1781__, new_new_n1782__, new_new_n1783__,
    new_new_n1784__, new_new_n1785__, new_new_n1786__, new_new_n1787__,
    new_new_n1788__, new_new_n1789__, new_new_n1790__, new_new_n1791__,
    new_new_n1792__, new_new_n1793__, new_new_n1794__, new_new_n1795__,
    new_new_n1796__, new_new_n1797__, new_new_n1798__, new_new_n1799__,
    new_new_n1800__, new_new_n1801__, new_new_n1802__, new_new_n1803__,
    new_new_n1804__, new_new_n1805__, new_new_n1806__, new_new_n1807__,
    new_new_n1808__, new_new_n1809__, new_new_n1810__, new_new_n1811__,
    new_new_n1812__, new_new_n1813__, new_new_n1814__, new_new_n1815__,
    new_new_n1816__, new_new_n1817__, new_new_n1818__, new_new_n1819__,
    new_new_n1820__, new_new_n1821__, new_new_n1822__, new_new_n1823__,
    new_new_n1824__, new_new_n1825__, new_new_n1826__, new_new_n1827__,
    new_new_n1828__, new_new_n1829__, new_new_n1830__, new_new_n1831__,
    new_new_n1832__, new_new_n1833__, new_new_n1834__, new_new_n1835__,
    new_new_n1836__, new_new_n1837__, new_new_n1838__, new_new_n1839__,
    new_new_n1840__, new_new_n1841__, new_new_n1842__, new_new_n1843__,
    new_new_n1844__, new_new_n1845__, new_new_n1846__, new_new_n1847__,
    new_new_n1848__, new_new_n1849__, new_new_n1850__, new_new_n1851__,
    new_new_n1852__, new_new_n1853__, new_new_n1854__, new_new_n1855__,
    new_new_n1856__, new_new_n1857__, new_new_n1858__, new_new_n1859__,
    new_new_n1860__, new_new_n1861__, new_new_n1862__, new_new_n1863__,
    new_new_n1864__, new_new_n1865__, new_new_n1866__, new_new_n1867__,
    new_new_n1868__, new_new_n1869__, new_new_n1870__, new_new_n1871__,
    new_new_n1872__, new_new_n1873__, new_new_n1874__, new_new_n1875__,
    new_new_n1876__, new_new_n1877__, new_new_n1878__, new_new_n1879__,
    new_new_n1880__, new_new_n1881__, new_new_n1882__, new_new_n1883__,
    new_new_n1884__, new_new_n1885__, new_new_n1886__, new_new_n1887__,
    new_new_n1888__, new_new_n1889__, new_new_n1890__, new_new_n1891__,
    new_new_n1892__, new_new_n1893__, new_new_n1894__, new_new_n1895__,
    new_new_n1896__, new_new_n1897__, new_new_n1898__, new_new_n1899__,
    new_new_n1900__, new_new_n1901__, new_new_n1902__, new_new_n1903__,
    new_new_n1904__, new_new_n1905__, new_new_n1906__, new_new_n1907__,
    new_new_n1908__, new_new_n1909__, new_new_n1910__, new_new_n1911__,
    new_new_n1912__, new_new_n1913__, new_new_n1914__, new_new_n1915__,
    new_new_n1916__, new_new_n1917__, new_new_n1918__, new_new_n1919__,
    new_new_n1920__, new_new_n1921__, new_new_n1922__, new_new_n1923__,
    new_new_n1924__, new_new_n1925__, new_new_n1926__, new_new_n1927__,
    new_new_n1928__, new_new_n1929__, new_new_n1930__, new_new_n1931__,
    new_new_n1932__, new_new_n1933__, new_new_n1934__, new_new_n1935__,
    new_new_n1936__, new_new_n1937__, new_new_n1938__, new_new_n1939__,
    new_new_n1940__, new_new_n1941__, new_new_n1942__, new_new_n1943__,
    new_new_n1944__, new_new_n1945__, new_new_n1946__, new_new_n1947__,
    new_new_n1948__, new_new_n1949__, new_new_n1950__, new_new_n1951__,
    new_new_n1952__, new_new_n1953__, new_new_n1954__, new_new_n1955__,
    new_new_n1956__, new_new_n1957__, new_new_n1958__, new_new_n1959__,
    new_new_n1960__, new_new_n1961__, new_new_n1962__, new_new_n1963__,
    new_new_n1964__, new_new_n1965__, new_new_n1966__, new_new_n1967__,
    new_new_n1968__, new_new_n1969__, new_new_n1970__, new_new_n1971__,
    new_new_n1972__, new_new_n1973__, new_new_n1974__, new_new_n1975__,
    new_new_n1976__, new_new_n1977__, new_new_n1978__, new_new_n1979__,
    new_new_n1980__, new_new_n1981__, new_new_n1982__, new_new_n1983__,
    new_new_n1984__, new_new_n1985__, new_new_n1986__, new_new_n1987__,
    new_new_n1988__, new_new_n1989__, new_new_n1990__, new_new_n1991__,
    new_new_n1992__, new_new_n1993__, new_new_n1994__, new_new_n1995__,
    new_new_n1996__, new_new_n1997__, new_new_n1998__, new_new_n1999__,
    new_new_n2000__, new_new_n2001__, new_new_n2002__, new_new_n2003__,
    new_new_n2004__, new_new_n2005__, new_new_n2006__, new_new_n2007__,
    new_new_n2008__, new_new_n2009__, new_new_n2010__, new_new_n2011__,
    new_new_n2012__, new_new_n2013__, new_new_n2014__, new_new_n2015__,
    new_new_n2016__, new_new_n2017__, new_new_n2018__, new_new_n2019__,
    new_new_n2020__, new_new_n2021__, new_new_n2022__, new_new_n2023__,
    new_new_n2024__, new_new_n2025__, new_new_n2026__, new_new_n2027__,
    new_new_n2028__, new_new_n2029__, new_new_n2030__, new_new_n2031__,
    new_new_n2032__, new_new_n2033__, new_new_n2034__, new_new_n2035__,
    new_new_n2036__, new_new_n2037__, new_new_n2038__, new_new_n2039__,
    new_new_n2040__, new_new_n2041__, new_new_n2042__, new_new_n2043__,
    new_new_n2044__, new_new_n2045__, new_new_n2046__, new_new_n2047__,
    new_new_n2048__, new_new_n2049__, new_new_n2050__, new_new_n2051__,
    new_new_n2052__, new_new_n2053__, new_new_n2054__, new_new_n2055__,
    new_new_n2056__, new_new_n2057__, new_new_n2058__, new_new_n2059__,
    new_new_n2060__, new_new_n2061__, new_new_n2062__, new_new_n2063__,
    new_new_n2064__, new_new_n2065__, new_new_n2066__, new_new_n2067__,
    new_new_n2068__, new_new_n2069__, new_new_n2070__, new_new_n2071__,
    new_new_n2072__, new_new_n2073__, new_new_n2074__, new_new_n2075__,
    new_new_n2076__, new_new_n2077__, new_new_n2078__, new_new_n2079__,
    new_new_n2080__, new_new_n2081__, new_new_n2082__, new_new_n2083__,
    new_new_n2084__, new_new_n2085__, new_new_n2086__, new_new_n2087__,
    new_new_n2088__, new_new_n2089__, new_new_n2090__, new_new_n2091__,
    new_new_n2092__, new_new_n2093__, new_new_n2094__, new_new_n2095__,
    new_new_n2096__, new_new_n2097__, new_new_n2098__, new_new_n2099__,
    new_new_n2100__, new_new_n2101__, new_new_n2102__, new_new_n2103__,
    new_new_n2104__, new_new_n2105__, new_new_n2106__, new_new_n2107__,
    new_new_n2108__, new_new_n2109__, new_new_n2110__, new_new_n2111__,
    new_new_n2112__, new_new_n2113__, new_new_n2114__, new_new_n2115__,
    new_new_n2116__, new_new_n2117__, new_new_n2118__, new_new_n2119__,
    new_new_n2120__, new_new_n2121__, new_new_n2122__, new_new_n2123__,
    new_new_n2124__, new_new_n2125__, new_new_n2126__, new_new_n2127__,
    new_new_n2128__, new_new_n2129__, new_new_n2130__, new_new_n2131__,
    new_new_n2132__, new_new_n2133__, new_new_n2134__, new_new_n2135__,
    new_new_n2136__, new_new_n2137__, new_new_n2138__, new_new_n2139__,
    new_new_n2140__, new_new_n2141__, new_new_n2142__, new_new_n2143__,
    new_new_n2144__, new_new_n2145__, new_new_n2146__, new_new_n2147__,
    new_new_n2148__, new_new_n2149__, new_new_n2150__, new_new_n2151__,
    new_new_n2152__, new_new_n2153__, new_new_n2154__, new_new_n2155__,
    new_new_n2156__, new_new_n2157__, new_new_n2158__, new_new_n2159__,
    new_new_n2160__, new_new_n2161__, new_new_n2162__, new_new_n2163__,
    new_new_n2164__, new_new_n2165__, new_new_n2166__, new_new_n2167__,
    new_new_n2168__, new_new_n2169__, new_new_n2170__, new_new_n2171__,
    new_new_n2172__, new_new_n2173__, new_new_n2174__, new_new_n2175__,
    new_new_n2176__, new_new_n2177__, new_new_n2178__, new_new_n2179__,
    new_new_n2180__, new_new_n2181__, new_new_n2182__, new_new_n2183__,
    new_new_n2184__, new_new_n2185__, new_new_n2186__, new_new_n2187__,
    new_new_n2188__, new_new_n2189__, new_new_n2190__, new_new_n2191__,
    new_new_n2192__, new_new_n2193__, new_new_n2194__, new_new_n2195__,
    new_new_n2196__, new_new_n2197__, new_new_n2198__, new_new_n2199__,
    new_new_n2200__, new_new_n2201__, new_new_n2202__, new_new_n2203__,
    new_new_n2204__, new_new_n2205__, new_new_n2206__, new_new_n2207__,
    new_new_n2208__, new_new_n2209__, new_new_n2210__, new_new_n2211__,
    new_new_n2212__, new_new_n2213__, new_new_n2214__, new_new_n2215__,
    new_new_n2216__, new_new_n2217__, new_new_n2218__, new_new_n2219__,
    new_new_n2220__, new_new_n2221__, new_new_n2222__, new_new_n2223__,
    new_new_n2224__, new_new_n2225__, new_new_n2226__, new_new_n2227__,
    new_new_n2228__, new_new_n2229__, new_new_n2230__, new_new_n2231__,
    new_new_n2232__, new_new_n2233__, new_new_n2234__, new_new_n2235__,
    new_new_n2236__, new_new_n2237__, new_new_n2238__, new_new_n2239__,
    new_new_n2240__, new_new_n2241__, new_new_n2242__, new_new_n2243__,
    new_new_n2244__, new_new_n2245__, new_new_n2246__, new_new_n2247__,
    new_new_n2248__, new_new_n2249__, new_new_n2250__, new_new_n2251__,
    new_new_n2252__, new_new_n2253__, new_new_n2254__, new_new_n2255__,
    new_new_n2256__, new_new_n2257__, new_new_n2258__, new_new_n2259__,
    new_new_n2260__, new_new_n2261__, new_new_n2262__, new_new_n2263__,
    new_new_n2264__, new_new_n2265__, new_new_n2266__, new_new_n2267__,
    new_new_n2268__, new_new_n2269__, new_new_n2270__, new_new_n2271__,
    new_new_n2272__, new_new_n2273__, new_new_n2274__, new_new_n2275__,
    n3791, n3794, n3797, n3800, n3803, n3806, n3809, n3812, n3815, n3818,
    n3821, n3824, n3827, n3830, n3833, n3836, n3839, n3842, n3845, n3848,
    n3851, n3854, n3857, n3860, n3863, n3866, n3869, n3872, n3875, n3878,
    n3881, n3884, n3887, n3890, n3893, n3896, n3899, n3902, n3905, n3908,
    n3911, n3914, n3917, n3920, n3923, n3926, n3929, n3932, n3935, n3938,
    n3941, n3944, n3947, n3950, n3953, n3956, n3959, n3962, n3965, n3968,
    n3971, n3974, n3977, n3980, n3983, n3986, n3989, n3992, n3995, n3998,
    n4001, n4004, n4007, n4010, n4013, n4016, n4019, n4022, n4025, n4028,
    n4031, n4034, n4037, n4040, n4043, n4046, n4049, n4052, n4055, n4058,
    n4061, n4064, n4067, n4070, n4073, n4076, n4079, n4082, n4085, n4088,
    n4091, n4094, n4097, n4100, n4103, n4106, n4109, n4112, n4115, n4118,
    n4121, n4124, n4127, n4130, n4133, n4136, n4139, n4142, n4145, n4148,
    n4151, n4154, n4157, n4160, n4163, n4166, n4169, n4172, n4175, n4178,
    n4181, n4184, n4187, n4190, n4193, n4196, n4199, n4202, n4205, n4208,
    n4211, n4214, n4217, n4220, n4223, n4226, n4229, n4232, n4235, n4238,
    n4241, n4244, n4247, n4250, n4253, n4256, n4259, n4262, n4265, n4268,
    n4271, n4274, n4277, n4280, n4283, n4286, n4289, n4292, n4295, n4298,
    n4301, n4304, n4307, n4310, n4313, n4316, n4319, n4322, n4325, n4328,
    n4331, n4334, n4337, n4340, n4343, n4346, n4349, n4352;
  not1  g0000(.din(G1), .dout(new_new_n451__));
  not1  g0001(.din(G2), .dout(new_new_n453__));
  not1  g0002(.din(G3), .dout(new_new_n455__));
  not1  g0003(.din(G4), .dout(new_new_n457__));
  not1  g0004(.din(G5), .dout(new_new_n459__));
  not1  g0005(.din(G6), .dout(new_new_n461__));
  not1  g0006(.din(G7), .dout(new_new_n463__));
  not1  g0007(.din(G8), .dout(new_new_n465__));
  not1  g0008(.din(G9), .dout(new_new_n467__));
  not1  g0009(.din(G10), .dout(new_new_n469__));
  not1  g0010(.din(G11), .dout(new_new_n471__));
  not1  g0011(.din(G12), .dout(new_new_n473__));
  not1  g0012(.din(G13), .dout(new_new_n475__));
  not1  g0013(.din(G14), .dout(new_new_n477__));
  not1  g0014(.din(G15), .dout(new_new_n479__));
  not1  g0015(.din(G16), .dout(new_new_n481__));
  not1  g0016(.din(G17), .dout(new_new_n483__));
  not1  g0017(.din(G18), .dout(new_new_n485__));
  not1  g0018(.din(G19), .dout(new_new_n487__));
  not1  g0019(.din(G20), .dout(new_new_n489__));
  not1  g0020(.din(G21), .dout(new_new_n491__));
  not1  g0021(.din(G22), .dout(new_new_n493__));
  not1  g0022(.din(G23), .dout(new_new_n495__));
  not1  g0023(.din(G24), .dout(new_new_n497__));
  not1  g0024(.din(G25), .dout(new_new_n499__));
  not1  g0025(.din(G26), .dout(new_new_n501__));
  not1  g0026(.din(G27), .dout(new_new_n503__));
  not1  g0027(.din(G28), .dout(new_new_n505__));
  not1  g0028(.din(G29), .dout(new_new_n507__));
  not1  g0029(.din(G30), .dout(new_new_n509__));
  not1  g0030(.din(G31), .dout(new_new_n511__));
  not1  g0031(.din(G32), .dout(new_new_n513__));
  not1  g0032(.din(G33), .dout(new_new_n515__));
  not1  g0033(.din(G34), .dout(new_new_n517__));
  not1  g0034(.din(G35), .dout(new_new_n519__));
  not1  g0035(.din(G36), .dout(new_new_n521__));
  not1  g0036(.din(G37), .dout(new_new_n523__));
  not1  g0037(.din(G38), .dout(new_new_n525__));
  not1  g0038(.din(G39), .dout(new_new_n527__));
  not1  g0039(.din(G40), .dout(new_new_n529__));
  not1  g0040(.din(G41), .dout(new_new_n531__));
  buf1  g0041(.din(n286_lo), .dout(new_new_n532__));
  not1  g0042(.din(n286_lo), .dout(new_new_n533__));
  buf1  g0043(.din(n298_lo), .dout(new_new_n534__));
  not1  g0044(.din(n298_lo), .dout(new_new_n535__));
  buf1  g0045(.din(n310_lo), .dout(new_new_n536__));
  not1  g0046(.din(n310_lo), .dout(new_new_n537__));
  buf1  g0047(.din(n322_lo), .dout(new_new_n538__));
  not1  g0048(.din(n322_lo), .dout(new_new_n539__));
  buf1  g0049(.din(n334_lo), .dout(new_new_n540__));
  not1  g0050(.din(n334_lo), .dout(new_new_n541__));
  buf1  g0051(.din(n346_lo), .dout(new_new_n542__));
  not1  g0052(.din(n346_lo), .dout(new_new_n543__));
  buf1  g0053(.din(n358_lo), .dout(new_new_n544__));
  not1  g0054(.din(n358_lo), .dout(new_new_n545__));
  buf1  g0055(.din(n370_lo), .dout(new_new_n546__));
  not1  g0056(.din(n370_lo), .dout(new_new_n547__));
  buf1  g0057(.din(n382_lo), .dout(new_new_n548__));
  not1  g0058(.din(n382_lo), .dout(new_new_n549__));
  buf1  g0059(.din(n394_lo), .dout(new_new_n550__));
  not1  g0060(.din(n394_lo), .dout(new_new_n551__));
  buf1  g0061(.din(n406_lo), .dout(new_new_n552__));
  not1  g0062(.din(n406_lo), .dout(new_new_n553__));
  buf1  g0063(.din(n418_lo), .dout(new_new_n554__));
  not1  g0064(.din(n418_lo), .dout(new_new_n555__));
  buf1  g0065(.din(n430_lo), .dout(new_new_n556__));
  not1  g0066(.din(n430_lo), .dout(new_new_n557__));
  buf1  g0067(.din(n442_lo), .dout(new_new_n558__));
  not1  g0068(.din(n442_lo), .dout(new_new_n559__));
  buf1  g0069(.din(n454_lo), .dout(new_new_n560__));
  not1  g0070(.din(n454_lo), .dout(new_new_n561__));
  buf1  g0071(.din(n466_lo), .dout(new_new_n562__));
  not1  g0072(.din(n466_lo), .dout(new_new_n563__));
  buf1  g0073(.din(n478_lo), .dout(new_new_n564__));
  not1  g0074(.din(n478_lo), .dout(new_new_n565__));
  buf1  g0075(.din(n490_lo), .dout(new_new_n566__));
  not1  g0076(.din(n490_lo), .dout(new_new_n567__));
  buf1  g0077(.din(n502_lo), .dout(new_new_n568__));
  not1  g0078(.din(n502_lo), .dout(new_new_n569__));
  buf1  g0079(.din(n514_lo), .dout(new_new_n570__));
  not1  g0080(.din(n514_lo), .dout(new_new_n571__));
  buf1  g0081(.din(n526_lo), .dout(new_new_n572__));
  not1  g0082(.din(n526_lo), .dout(new_new_n573__));
  buf1  g0083(.din(n538_lo), .dout(new_new_n574__));
  not1  g0084(.din(n538_lo), .dout(new_new_n575__));
  buf1  g0085(.din(n550_lo), .dout(new_new_n576__));
  not1  g0086(.din(n550_lo), .dout(new_new_n577__));
  buf1  g0087(.din(n562_lo), .dout(new_new_n578__));
  not1  g0088(.din(n562_lo), .dout(new_new_n579__));
  buf1  g0089(.din(n574_lo), .dout(new_new_n580__));
  not1  g0090(.din(n574_lo), .dout(new_new_n581__));
  buf1  g0091(.din(n586_lo), .dout(new_new_n582__));
  not1  g0092(.din(n586_lo), .dout(new_new_n583__));
  buf1  g0093(.din(n598_lo), .dout(new_new_n584__));
  not1  g0094(.din(n598_lo), .dout(new_new_n585__));
  buf1  g0095(.din(n610_lo), .dout(new_new_n586__));
  not1  g0096(.din(n610_lo), .dout(new_new_n587__));
  buf1  g0097(.din(n622_lo), .dout(new_new_n588__));
  not1  g0098(.din(n622_lo), .dout(new_new_n589__));
  buf1  g0099(.din(n634_lo), .dout(new_new_n590__));
  not1  g0100(.din(n634_lo), .dout(new_new_n591__));
  buf1  g0101(.din(n646_lo), .dout(new_new_n592__));
  not1  g0102(.din(n646_lo), .dout(new_new_n593__));
  buf1  g0103(.din(n658_lo), .dout(new_new_n594__));
  not1  g0104(.din(n658_lo), .dout(new_new_n595__));
  not1  g0105(.din(n661_lo), .dout(new_new_n597__));
  not1  g0106(.din(n673_lo), .dout(new_new_n599__));
  not1  g0107(.din(n685_lo), .dout(new_new_n601__));
  not1  g0108(.din(n697_lo), .dout(new_new_n603__));
  not1  g0109(.din(n709_lo), .dout(new_new_n605__));
  not1  g0110(.din(n721_lo), .dout(new_new_n607__));
  not1  g0111(.din(n733_lo), .dout(new_new_n609__));
  not1  g0112(.din(n745_lo), .dout(new_new_n611__));
  not1  g0113(.din(n757_lo), .dout(new_new_n613__));
  buf1  g0114(.din(n1248_o2), .dout(new_new_n614__));
  not1  g0115(.din(n1248_o2), .dout(new_new_n615__));
  buf1  g0116(.din(n1249_o2), .dout(new_new_n616__));
  not1  g0117(.din(n1249_o2), .dout(new_new_n617__));
  buf1  g0118(.din(n1250_o2), .dout(new_new_n618__));
  not1  g0119(.din(n1250_o2), .dout(new_new_n619__));
  buf1  g0120(.din(n1251_o2), .dout(new_new_n620__));
  not1  g0121(.din(n1251_o2), .dout(new_new_n621__));
  buf1  g0122(.din(n1252_o2), .dout(new_new_n622__));
  not1  g0123(.din(n1252_o2), .dout(new_new_n623__));
  buf1  g0124(.din(n1253_o2), .dout(new_new_n624__));
  not1  g0125(.din(n1253_o2), .dout(new_new_n625__));
  buf1  g0126(.din(n1254_o2), .dout(new_new_n626__));
  not1  g0127(.din(n1254_o2), .dout(new_new_n627__));
  buf1  g0128(.din(n1255_o2), .dout(new_new_n628__));
  not1  g0129(.din(n1255_o2), .dout(new_new_n629__));
  not1  g0130(.din(n1207_o2), .dout(new_new_n631__));
  not1  g0131(.din(n1208_o2), .dout(new_new_n633__));
  not1  g0132(.din(n1209_o2), .dout(new_new_n635__));
  not1  g0133(.din(n1210_o2), .dout(new_new_n637__));
  not1  g0134(.din(n1211_o2), .dout(new_new_n639__));
  not1  g0135(.din(n1212_o2), .dout(new_new_n641__));
  not1  g0136(.din(n1213_o2), .dout(new_new_n643__));
  not1  g0137(.din(n1214_o2), .dout(new_new_n645__));
  not1  g0138(.din(n1215_o2), .dout(new_new_n647__));
  not1  g0139(.din(n1216_o2), .dout(new_new_n649__));
  not1  g0140(.din(n1217_o2), .dout(new_new_n651__));
  not1  g0141(.din(n1218_o2), .dout(new_new_n653__));
  not1  g0142(.din(n1219_o2), .dout(new_new_n655__));
  not1  g0143(.din(n1220_o2), .dout(new_new_n657__));
  not1  g0144(.din(n1221_o2), .dout(new_new_n659__));
  not1  g0145(.din(n1222_o2), .dout(new_new_n661__));
  not1  g0146(.din(n1223_o2), .dout(new_new_n663__));
  not1  g0147(.din(n1224_o2), .dout(new_new_n665__));
  not1  g0148(.din(n1225_o2), .dout(new_new_n667__));
  not1  g0149(.din(n1226_o2), .dout(new_new_n669__));
  not1  g0150(.din(n1227_o2), .dout(new_new_n671__));
  not1  g0151(.din(n1228_o2), .dout(new_new_n673__));
  not1  g0152(.din(n1229_o2), .dout(new_new_n675__));
  not1  g0153(.din(n1230_o2), .dout(new_new_n677__));
  not1  g0154(.din(n1231_o2), .dout(new_new_n679__));
  not1  g0155(.din(n1232_o2), .dout(new_new_n681__));
  not1  g0156(.din(n1233_o2), .dout(new_new_n683__));
  not1  g0157(.din(n1234_o2), .dout(new_new_n685__));
  not1  g0158(.din(n1235_o2), .dout(new_new_n687__));
  not1  g0159(.din(n1236_o2), .dout(new_new_n689__));
  not1  g0160(.din(n1237_o2), .dout(new_new_n691__));
  not1  g0161(.din(n1238_o2), .dout(new_new_n693__));
  buf1  g0162(.din(G374_o2), .dout(new_new_n694__));
  not1  g0163(.din(G374_o2), .dout(new_new_n695__));
  buf1  g0164(.din(G376_o2), .dout(new_new_n696__));
  not1  g0165(.din(G376_o2), .dout(new_new_n697__));
  buf1  g0166(.din(G370_o2), .dout(new_new_n698__));
  not1  g0167(.din(G370_o2), .dout(new_new_n699__));
  buf1  g0168(.din(G372_o2), .dout(new_new_n700__));
  not1  g0169(.din(G372_o2), .dout(new_new_n701__));
  buf1  g0170(.din(G373_o2), .dout(new_new_n702__));
  not1  g0171(.din(G373_o2), .dout(new_new_n703__));
  buf1  g0172(.din(G377_o2), .dout(new_new_n704__));
  not1  g0173(.din(G377_o2), .dout(new_new_n705__));
  buf1  g0174(.din(G371_o2), .dout(new_new_n706__));
  not1  g0175(.din(G371_o2), .dout(new_new_n707__));
  buf1  g0176(.din(G375_o2), .dout(new_new_n708__));
  not1  g0177(.din(G375_o2), .dout(new_new_n709__));
  buf1  g0178(.din(G354_o2), .dout(new_new_n710__));
  not1  g0179(.din(G354_o2), .dout(new_new_n711__));
  buf1  g0180(.din(G356_o2), .dout(new_new_n712__));
  not1  g0181(.din(G356_o2), .dout(new_new_n713__));
  buf1  g0182(.din(G350_o2), .dout(new_new_n714__));
  not1  g0183(.din(G350_o2), .dout(new_new_n715__));
  buf1  g0184(.din(G352_o2), .dout(new_new_n716__));
  not1  g0185(.din(G352_o2), .dout(new_new_n717__));
  buf1  g0186(.din(G353_o2), .dout(new_new_n718__));
  not1  g0187(.din(G353_o2), .dout(new_new_n719__));
  buf1  g0188(.din(G357_o2), .dout(new_new_n720__));
  not1  g0189(.din(G357_o2), .dout(new_new_n721__));
  buf1  g0190(.din(G351_o2), .dout(new_new_n722__));
  not1  g0191(.din(G351_o2), .dout(new_new_n723__));
  buf1  g0192(.din(G355_o2), .dout(new_new_n724__));
  not1  g0193(.din(G355_o2), .dout(new_new_n725__));
  buf1  g0194(.din(G386_o2), .dout(new_new_n726__));
  not1  g0195(.din(G386_o2), .dout(new_new_n727__));
  buf1  g0196(.din(G391_o2), .dout(new_new_n728__));
  not1  g0197(.din(G391_o2), .dout(new_new_n729__));
  buf1  g0198(.din(n283_lo_buf_o2), .dout(new_new_n730__));
  not1  g0199(.din(n283_lo_buf_o2), .dout(new_new_n731__));
  buf1  g0200(.din(n295_lo_buf_o2), .dout(new_new_n732__));
  not1  g0201(.din(n295_lo_buf_o2), .dout(new_new_n733__));
  buf1  g0202(.din(n307_lo_buf_o2), .dout(new_new_n734__));
  not1  g0203(.din(n307_lo_buf_o2), .dout(new_new_n735__));
  buf1  g0204(.din(n319_lo_buf_o2), .dout(new_new_n736__));
  not1  g0205(.din(n319_lo_buf_o2), .dout(new_new_n737__));
  buf1  g0206(.din(n331_lo_buf_o2), .dout(new_new_n738__));
  not1  g0207(.din(n331_lo_buf_o2), .dout(new_new_n739__));
  buf1  g0208(.din(n343_lo_buf_o2), .dout(new_new_n740__));
  not1  g0209(.din(n343_lo_buf_o2), .dout(new_new_n741__));
  buf1  g0210(.din(n355_lo_buf_o2), .dout(new_new_n742__));
  not1  g0211(.din(n355_lo_buf_o2), .dout(new_new_n743__));
  buf1  g0212(.din(n367_lo_buf_o2), .dout(new_new_n744__));
  not1  g0213(.din(n367_lo_buf_o2), .dout(new_new_n745__));
  buf1  g0214(.din(n379_lo_buf_o2), .dout(new_new_n746__));
  not1  g0215(.din(n379_lo_buf_o2), .dout(new_new_n747__));
  buf1  g0216(.din(n391_lo_buf_o2), .dout(new_new_n748__));
  not1  g0217(.din(n391_lo_buf_o2), .dout(new_new_n749__));
  buf1  g0218(.din(n403_lo_buf_o2), .dout(new_new_n750__));
  not1  g0219(.din(n403_lo_buf_o2), .dout(new_new_n751__));
  buf1  g0220(.din(n415_lo_buf_o2), .dout(new_new_n752__));
  not1  g0221(.din(n415_lo_buf_o2), .dout(new_new_n753__));
  buf1  g0222(.din(n427_lo_buf_o2), .dout(new_new_n754__));
  not1  g0223(.din(n427_lo_buf_o2), .dout(new_new_n755__));
  buf1  g0224(.din(n439_lo_buf_o2), .dout(new_new_n756__));
  not1  g0225(.din(n439_lo_buf_o2), .dout(new_new_n757__));
  buf1  g0226(.din(n451_lo_buf_o2), .dout(new_new_n758__));
  not1  g0227(.din(n451_lo_buf_o2), .dout(new_new_n759__));
  buf1  g0228(.din(n463_lo_buf_o2), .dout(new_new_n760__));
  not1  g0229(.din(n463_lo_buf_o2), .dout(new_new_n761__));
  buf1  g0230(.din(n475_lo_buf_o2), .dout(new_new_n762__));
  not1  g0231(.din(n475_lo_buf_o2), .dout(new_new_n763__));
  buf1  g0232(.din(n487_lo_buf_o2), .dout(new_new_n764__));
  not1  g0233(.din(n487_lo_buf_o2), .dout(new_new_n765__));
  buf1  g0234(.din(n499_lo_buf_o2), .dout(new_new_n766__));
  not1  g0235(.din(n499_lo_buf_o2), .dout(new_new_n767__));
  buf1  g0236(.din(n511_lo_buf_o2), .dout(new_new_n768__));
  not1  g0237(.din(n511_lo_buf_o2), .dout(new_new_n769__));
  buf1  g0238(.din(n523_lo_buf_o2), .dout(new_new_n770__));
  not1  g0239(.din(n523_lo_buf_o2), .dout(new_new_n771__));
  buf1  g0240(.din(n535_lo_buf_o2), .dout(new_new_n772__));
  not1  g0241(.din(n535_lo_buf_o2), .dout(new_new_n773__));
  buf1  g0242(.din(n547_lo_buf_o2), .dout(new_new_n774__));
  not1  g0243(.din(n547_lo_buf_o2), .dout(new_new_n775__));
  buf1  g0244(.din(n559_lo_buf_o2), .dout(new_new_n776__));
  not1  g0245(.din(n559_lo_buf_o2), .dout(new_new_n777__));
  buf1  g0246(.din(n571_lo_buf_o2), .dout(new_new_n778__));
  not1  g0247(.din(n571_lo_buf_o2), .dout(new_new_n779__));
  buf1  g0248(.din(n583_lo_buf_o2), .dout(new_new_n780__));
  not1  g0249(.din(n583_lo_buf_o2), .dout(new_new_n781__));
  buf1  g0250(.din(n595_lo_buf_o2), .dout(new_new_n782__));
  not1  g0251(.din(n595_lo_buf_o2), .dout(new_new_n783__));
  buf1  g0252(.din(n607_lo_buf_o2), .dout(new_new_n784__));
  not1  g0253(.din(n607_lo_buf_o2), .dout(new_new_n785__));
  buf1  g0254(.din(n619_lo_buf_o2), .dout(new_new_n786__));
  not1  g0255(.din(n619_lo_buf_o2), .dout(new_new_n787__));
  buf1  g0256(.din(n631_lo_buf_o2), .dout(new_new_n788__));
  not1  g0257(.din(n631_lo_buf_o2), .dout(new_new_n789__));
  buf1  g0258(.din(n643_lo_buf_o2), .dout(new_new_n790__));
  not1  g0259(.din(n643_lo_buf_o2), .dout(new_new_n791__));
  buf1  g0260(.din(n655_lo_buf_o2), .dout(new_new_n792__));
  not1  g0261(.din(n655_lo_buf_o2), .dout(new_new_n793__));
  buf1  g0262(.din(G234_o2), .dout(new_new_n794__));
  not1  g0263(.din(G234_o2), .dout(new_new_n795__));
  buf1  g0264(.din(G247_o2), .dout(new_new_n796__));
  not1  g0265(.din(G247_o2), .dout(new_new_n797__));
  buf1  g0266(.din(G260_o2), .dout(new_new_n798__));
  not1  g0267(.din(G260_o2), .dout(new_new_n799__));
  buf1  g0268(.din(G273_o2), .dout(new_new_n800__));
  not1  g0269(.din(G273_o2), .dout(new_new_n801__));
  buf1  g0270(.din(G286_o2), .dout(new_new_n802__));
  not1  g0271(.din(G286_o2), .dout(new_new_n803__));
  buf1  g0272(.din(G299_o2), .dout(new_new_n804__));
  not1  g0273(.din(G299_o2), .dout(new_new_n805__));
  buf1  g0274(.din(G312_o2), .dout(new_new_n806__));
  not1  g0275(.din(G312_o2), .dout(new_new_n807__));
  buf1  g0276(.din(G325_o2), .dout(new_new_n808__));
  not1  g0277(.din(G325_o2), .dout(new_new_n809__));
  buf1  g0278(.din(n667_lo_buf_o2), .dout(new_new_n810__));
  not1  g0279(.din(n667_lo_buf_o2), .dout(new_new_n811__));
  buf1  g0280(.din(n679_lo_buf_o2), .dout(new_new_n812__));
  not1  g0281(.din(n679_lo_buf_o2), .dout(new_new_n813__));
  buf1  g0282(.din(n691_lo_buf_o2), .dout(new_new_n814__));
  not1  g0283(.din(n691_lo_buf_o2), .dout(new_new_n815__));
  buf1  g0284(.din(n703_lo_buf_o2), .dout(new_new_n816__));
  not1  g0285(.din(n703_lo_buf_o2), .dout(new_new_n817__));
  buf1  g0286(.din(n715_lo_buf_o2), .dout(new_new_n818__));
  not1  g0287(.din(n715_lo_buf_o2), .dout(new_new_n819__));
  buf1  g0288(.din(n727_lo_buf_o2), .dout(new_new_n820__));
  not1  g0289(.din(n727_lo_buf_o2), .dout(new_new_n821__));
  buf1  g0290(.din(n739_lo_buf_o2), .dout(new_new_n822__));
  not1  g0291(.din(n739_lo_buf_o2), .dout(new_new_n823__));
  buf1  g0292(.din(n751_lo_buf_o2), .dout(new_new_n824__));
  not1  g0293(.din(n751_lo_buf_o2), .dout(new_new_n825__));
  buf1  g0294(.din(n763_lo_buf_o2), .dout(new_new_n826__));
  not1  g0295(.din(n763_lo_buf_o2), .dout(new_new_n827__));
  buf1  g0296(.din(G186_o2), .dout(new_new_n828__));
  not1  g0297(.din(G186_o2), .dout(new_new_n829__));
  buf1  g0298(.din(G189_o2), .dout(new_new_n830__));
  not1  g0299(.din(G189_o2), .dout(new_new_n831__));
  buf1  g0300(.din(G192_o2), .dout(new_new_n832__));
  not1  g0301(.din(G192_o2), .dout(new_new_n833__));
  buf1  g0302(.din(G195_o2), .dout(new_new_n834__));
  not1  g0303(.din(G195_o2), .dout(new_new_n835__));
  buf1  g0304(.din(G198_o2), .dout(new_new_n836__));
  not1  g0305(.din(G198_o2), .dout(new_new_n837__));
  buf1  g0306(.din(G201_o2), .dout(new_new_n838__));
  not1  g0307(.din(G201_o2), .dout(new_new_n839__));
  buf1  g0308(.din(G204_o2), .dout(new_new_n840__));
  not1  g0309(.din(G204_o2), .dout(new_new_n841__));
  buf1  g0310(.din(G207_o2), .dout(new_new_n842__));
  not1  g0311(.din(G207_o2), .dout(new_new_n843__));
  buf1  g0312(.din(n280_lo_buf_o2), .dout(new_new_n844__));
  not1  g0313(.din(n280_lo_buf_o2), .dout(new_new_n845__));
  buf1  g0314(.din(n292_lo_buf_o2), .dout(new_new_n846__));
  not1  g0315(.din(n292_lo_buf_o2), .dout(new_new_n847__));
  buf1  g0316(.din(n304_lo_buf_o2), .dout(new_new_n848__));
  not1  g0317(.din(n304_lo_buf_o2), .dout(new_new_n849__));
  buf1  g0318(.din(n316_lo_buf_o2), .dout(new_new_n850__));
  not1  g0319(.din(n316_lo_buf_o2), .dout(new_new_n851__));
  buf1  g0320(.din(n328_lo_buf_o2), .dout(new_new_n852__));
  not1  g0321(.din(n328_lo_buf_o2), .dout(new_new_n853__));
  buf1  g0322(.din(n340_lo_buf_o2), .dout(new_new_n854__));
  not1  g0323(.din(n340_lo_buf_o2), .dout(new_new_n855__));
  buf1  g0324(.din(n352_lo_buf_o2), .dout(new_new_n856__));
  not1  g0325(.din(n352_lo_buf_o2), .dout(new_new_n857__));
  buf1  g0326(.din(n364_lo_buf_o2), .dout(new_new_n858__));
  not1  g0327(.din(n364_lo_buf_o2), .dout(new_new_n859__));
  buf1  g0328(.din(n376_lo_buf_o2), .dout(new_new_n860__));
  not1  g0329(.din(n376_lo_buf_o2), .dout(new_new_n861__));
  buf1  g0330(.din(n388_lo_buf_o2), .dout(new_new_n862__));
  not1  g0331(.din(n388_lo_buf_o2), .dout(new_new_n863__));
  buf1  g0332(.din(n400_lo_buf_o2), .dout(new_new_n864__));
  not1  g0333(.din(n400_lo_buf_o2), .dout(new_new_n865__));
  buf1  g0334(.din(n412_lo_buf_o2), .dout(new_new_n866__));
  not1  g0335(.din(n412_lo_buf_o2), .dout(new_new_n867__));
  buf1  g0336(.din(n424_lo_buf_o2), .dout(new_new_n868__));
  not1  g0337(.din(n424_lo_buf_o2), .dout(new_new_n869__));
  buf1  g0338(.din(n436_lo_buf_o2), .dout(new_new_n870__));
  not1  g0339(.din(n436_lo_buf_o2), .dout(new_new_n871__));
  buf1  g0340(.din(n448_lo_buf_o2), .dout(new_new_n872__));
  not1  g0341(.din(n448_lo_buf_o2), .dout(new_new_n873__));
  buf1  g0342(.din(n460_lo_buf_o2), .dout(new_new_n874__));
  not1  g0343(.din(n460_lo_buf_o2), .dout(new_new_n875__));
  buf1  g0344(.din(n472_lo_buf_o2), .dout(new_new_n876__));
  not1  g0345(.din(n472_lo_buf_o2), .dout(new_new_n877__));
  buf1  g0346(.din(n484_lo_buf_o2), .dout(new_new_n878__));
  not1  g0347(.din(n484_lo_buf_o2), .dout(new_new_n879__));
  buf1  g0348(.din(n496_lo_buf_o2), .dout(new_new_n880__));
  not1  g0349(.din(n496_lo_buf_o2), .dout(new_new_n881__));
  buf1  g0350(.din(n508_lo_buf_o2), .dout(new_new_n882__));
  not1  g0351(.din(n508_lo_buf_o2), .dout(new_new_n883__));
  buf1  g0352(.din(n520_lo_buf_o2), .dout(new_new_n884__));
  not1  g0353(.din(n520_lo_buf_o2), .dout(new_new_n885__));
  buf1  g0354(.din(n532_lo_buf_o2), .dout(new_new_n886__));
  not1  g0355(.din(n532_lo_buf_o2), .dout(new_new_n887__));
  buf1  g0356(.din(n544_lo_buf_o2), .dout(new_new_n888__));
  not1  g0357(.din(n544_lo_buf_o2), .dout(new_new_n889__));
  buf1  g0358(.din(n556_lo_buf_o2), .dout(new_new_n890__));
  not1  g0359(.din(n556_lo_buf_o2), .dout(new_new_n891__));
  buf1  g0360(.din(n568_lo_buf_o2), .dout(new_new_n892__));
  not1  g0361(.din(n568_lo_buf_o2), .dout(new_new_n893__));
  buf1  g0362(.din(n580_lo_buf_o2), .dout(new_new_n894__));
  not1  g0363(.din(n580_lo_buf_o2), .dout(new_new_n895__));
  buf1  g0364(.din(n592_lo_buf_o2), .dout(new_new_n896__));
  not1  g0365(.din(n592_lo_buf_o2), .dout(new_new_n897__));
  buf1  g0366(.din(n604_lo_buf_o2), .dout(new_new_n898__));
  not1  g0367(.din(n604_lo_buf_o2), .dout(new_new_n899__));
  buf1  g0368(.din(n616_lo_buf_o2), .dout(new_new_n900__));
  not1  g0369(.din(n616_lo_buf_o2), .dout(new_new_n901__));
  buf1  g0370(.din(n628_lo_buf_o2), .dout(new_new_n902__));
  not1  g0371(.din(n628_lo_buf_o2), .dout(new_new_n903__));
  buf1  g0372(.din(n640_lo_buf_o2), .dout(new_new_n904__));
  not1  g0373(.din(n640_lo_buf_o2), .dout(new_new_n905__));
  buf1  g0374(.din(n652_lo_buf_o2), .dout(new_new_n906__));
  not1  g0375(.din(n652_lo_buf_o2), .dout(new_new_n907__));
  and1  g0376(.dina(new_new_n715__), .dinb(new_new_n1782__), .dout(new_new_n908__));
  or1   g0377(.dina(new_new_n714__), .dinb(new_new_n1787__), .dout(new_new_n909__));
  and1  g0378(.dina(new_new_n908__), .dinb(new_new_n1792__), .dout(new_new_n910__));
  or1   g0379(.dina(new_new_n909__), .dinb(new_new_n1797__), .dout(new_new_n911__));
  and1  g0380(.dina(new_new_n910__), .dinb(new_new_n723__), .dout(new_new_n912__));
  or1   g0381(.dina(new_new_n911__), .dinb(new_new_n722__), .dout(new_new_n913__));
  and1  g0382(.dina(new_new_n912__), .dinb(new_new_n1801__), .dout(new_new_n914__));
  or1   g0383(.dina(new_new_n913__), .dinb(new_new_n1804__), .dout(new_new_n915__));
  and1  g0384(.dina(new_new_n1807__), .dinb(new_new_n1811__), .dout(new_new_n916__));
  or1   g0385(.dina(new_new_n1815__), .dinb(new_new_n1819__), .dout(new_new_n917__));
  or1   g0386(.dina(new_new_n917__), .dinb(new_new_n532__), .dout(new_new_n918__));
  or1   g0387(.dina(new_new_n916__), .dinb(new_new_n533__), .dout(new_new_n919__));
  and1  g0388(.dina(new_new_n919__), .dinb(new_new_n918__), .dout(new_new_n920__));
  and1  g0389(.dina(new_new_n1807__), .dinb(new_new_n1824__), .dout(new_new_n921__));
  or1   g0390(.dina(new_new_n1815__), .dinb(new_new_n1829__), .dout(new_new_n922__));
  or1   g0391(.dina(new_new_n922__), .dinb(new_new_n534__), .dout(new_new_n923__));
  or1   g0392(.dina(new_new_n921__), .dinb(new_new_n535__), .dout(new_new_n924__));
  and1  g0393(.dina(new_new_n924__), .dinb(new_new_n923__), .dout(new_new_n925__));
  and1  g0394(.dina(new_new_n1808__), .dinb(new_new_n1834__), .dout(new_new_n926__));
  or1   g0395(.dina(new_new_n1816__), .dinb(new_new_n1839__), .dout(new_new_n927__));
  or1   g0396(.dina(new_new_n927__), .dinb(new_new_n536__), .dout(new_new_n928__));
  or1   g0397(.dina(new_new_n926__), .dinb(new_new_n537__), .dout(new_new_n929__));
  and1  g0398(.dina(new_new_n929__), .dinb(new_new_n928__), .dout(new_new_n930__));
  and1  g0399(.dina(new_new_n1808__), .dinb(new_new_n1844__), .dout(new_new_n931__));
  or1   g0400(.dina(new_new_n1816__), .dinb(new_new_n1849__), .dout(new_new_n932__));
  or1   g0401(.dina(new_new_n932__), .dinb(new_new_n538__), .dout(new_new_n933__));
  or1   g0402(.dina(new_new_n931__), .dinb(new_new_n539__), .dout(new_new_n934__));
  and1  g0403(.dina(new_new_n934__), .dinb(new_new_n933__), .dout(new_new_n935__));
  and1  g0404(.dina(new_new_n717__), .dinb(new_new_n1782__), .dout(new_new_n936__));
  or1   g0405(.dina(new_new_n716__), .dinb(new_new_n1787__), .dout(new_new_n937__));
  and1  g0406(.dina(new_new_n936__), .dinb(new_new_n719__), .dout(new_new_n938__));
  or1   g0407(.dina(new_new_n937__), .dinb(new_new_n718__), .dout(new_new_n939__));
  and1  g0408(.dina(new_new_n938__), .dinb(new_new_n1854__), .dout(new_new_n940__));
  or1   g0409(.dina(new_new_n939__), .dinb(new_new_n1859__), .dout(new_new_n941__));
  and1  g0410(.dina(new_new_n940__), .dinb(new_new_n1801__), .dout(new_new_n942__));
  or1   g0411(.dina(new_new_n941__), .dinb(new_new_n1804__), .dout(new_new_n943__));
  and1  g0412(.dina(new_new_n1863__), .dinb(new_new_n1811__), .dout(new_new_n944__));
  or1   g0413(.dina(new_new_n1866__), .dinb(new_new_n1819__), .dout(new_new_n945__));
  or1   g0414(.dina(new_new_n945__), .dinb(new_new_n540__), .dout(new_new_n946__));
  or1   g0415(.dina(new_new_n944__), .dinb(new_new_n541__), .dout(new_new_n947__));
  and1  g0416(.dina(new_new_n947__), .dinb(new_new_n946__), .dout(new_new_n948__));
  and1  g0417(.dina(new_new_n1863__), .dinb(new_new_n1824__), .dout(new_new_n949__));
  or1   g0418(.dina(new_new_n1866__), .dinb(new_new_n1829__), .dout(new_new_n950__));
  or1   g0419(.dina(new_new_n950__), .dinb(new_new_n542__), .dout(new_new_n951__));
  or1   g0420(.dina(new_new_n949__), .dinb(new_new_n543__), .dout(new_new_n952__));
  and1  g0421(.dina(new_new_n952__), .dinb(new_new_n951__), .dout(new_new_n953__));
  and1  g0422(.dina(new_new_n1864__), .dinb(new_new_n1834__), .dout(new_new_n954__));
  or1   g0423(.dina(new_new_n1867__), .dinb(new_new_n1839__), .dout(new_new_n955__));
  or1   g0424(.dina(new_new_n955__), .dinb(new_new_n544__), .dout(new_new_n956__));
  or1   g0425(.dina(new_new_n954__), .dinb(new_new_n545__), .dout(new_new_n957__));
  and1  g0426(.dina(new_new_n957__), .dinb(new_new_n956__), .dout(new_new_n958__));
  and1  g0427(.dina(new_new_n1864__), .dinb(new_new_n1844__), .dout(new_new_n959__));
  or1   g0428(.dina(new_new_n1867__), .dinb(new_new_n1849__), .dout(new_new_n960__));
  or1   g0429(.dina(new_new_n960__), .dinb(new_new_n546__), .dout(new_new_n961__));
  or1   g0430(.dina(new_new_n959__), .dinb(new_new_n547__), .dout(new_new_n962__));
  and1  g0431(.dina(new_new_n962__), .dinb(new_new_n961__), .dout(new_new_n963__));
  and1  g0432(.dina(new_new_n711__), .dinb(new_new_n1870__), .dout(new_new_n964__));
  or1   g0433(.dina(new_new_n710__), .dinb(new_new_n1875__), .dout(new_new_n965__));
  and1  g0434(.dina(new_new_n964__), .dinb(new_new_n1792__), .dout(new_new_n966__));
  or1   g0435(.dina(new_new_n965__), .dinb(new_new_n1797__), .dout(new_new_n967__));
  and1  g0436(.dina(new_new_n966__), .dinb(new_new_n725__), .dout(new_new_n968__));
  or1   g0437(.dina(new_new_n967__), .dinb(new_new_n724__), .dout(new_new_n969__));
  and1  g0438(.dina(new_new_n968__), .dinb(new_new_n1802__), .dout(new_new_n970__));
  or1   g0439(.dina(new_new_n969__), .dinb(new_new_n1805__), .dout(new_new_n971__));
  and1  g0440(.dina(new_new_n1879__), .dinb(new_new_n1812__), .dout(new_new_n972__));
  or1   g0441(.dina(new_new_n1882__), .dinb(new_new_n1820__), .dout(new_new_n973__));
  or1   g0442(.dina(new_new_n973__), .dinb(new_new_n548__), .dout(new_new_n974__));
  or1   g0443(.dina(new_new_n972__), .dinb(new_new_n549__), .dout(new_new_n975__));
  and1  g0444(.dina(new_new_n975__), .dinb(new_new_n974__), .dout(new_new_n976__));
  and1  g0445(.dina(new_new_n1879__), .dinb(new_new_n1825__), .dout(new_new_n977__));
  or1   g0446(.dina(new_new_n1882__), .dinb(new_new_n1830__), .dout(new_new_n978__));
  or1   g0447(.dina(new_new_n978__), .dinb(new_new_n550__), .dout(new_new_n979__));
  or1   g0448(.dina(new_new_n977__), .dinb(new_new_n551__), .dout(new_new_n980__));
  and1  g0449(.dina(new_new_n980__), .dinb(new_new_n979__), .dout(new_new_n981__));
  and1  g0450(.dina(new_new_n1880__), .dinb(new_new_n1835__), .dout(new_new_n982__));
  or1   g0451(.dina(new_new_n1883__), .dinb(new_new_n1840__), .dout(new_new_n983__));
  or1   g0452(.dina(new_new_n983__), .dinb(new_new_n552__), .dout(new_new_n984__));
  or1   g0453(.dina(new_new_n982__), .dinb(new_new_n553__), .dout(new_new_n985__));
  and1  g0454(.dina(new_new_n985__), .dinb(new_new_n984__), .dout(new_new_n986__));
  and1  g0455(.dina(new_new_n1880__), .dinb(new_new_n1845__), .dout(new_new_n987__));
  or1   g0456(.dina(new_new_n1883__), .dinb(new_new_n1850__), .dout(new_new_n988__));
  or1   g0457(.dina(new_new_n988__), .dinb(new_new_n554__), .dout(new_new_n989__));
  or1   g0458(.dina(new_new_n987__), .dinb(new_new_n555__), .dout(new_new_n990__));
  and1  g0459(.dina(new_new_n990__), .dinb(new_new_n989__), .dout(new_new_n991__));
  and1  g0460(.dina(new_new_n713__), .dinb(new_new_n1870__), .dout(new_new_n992__));
  or1   g0461(.dina(new_new_n712__), .dinb(new_new_n1875__), .dout(new_new_n993__));
  and1  g0462(.dina(new_new_n992__), .dinb(new_new_n721__), .dout(new_new_n994__));
  or1   g0463(.dina(new_new_n993__), .dinb(new_new_n720__), .dout(new_new_n995__));
  and1  g0464(.dina(new_new_n994__), .dinb(new_new_n1854__), .dout(new_new_n996__));
  or1   g0465(.dina(new_new_n995__), .dinb(new_new_n1859__), .dout(new_new_n997__));
  and1  g0466(.dina(new_new_n996__), .dinb(new_new_n1802__), .dout(new_new_n998__));
  or1   g0467(.dina(new_new_n997__), .dinb(new_new_n1805__), .dout(new_new_n999__));
  and1  g0468(.dina(new_new_n1885__), .dinb(new_new_n1812__), .dout(new_new_n1000__));
  or1   g0469(.dina(new_new_n1888__), .dinb(new_new_n1820__), .dout(new_new_n1001__));
  or1   g0470(.dina(new_new_n1001__), .dinb(new_new_n556__), .dout(new_new_n1002__));
  or1   g0471(.dina(new_new_n1000__), .dinb(new_new_n557__), .dout(new_new_n1003__));
  and1  g0472(.dina(new_new_n1003__), .dinb(new_new_n1002__), .dout(new_new_n1004__));
  and1  g0473(.dina(new_new_n1885__), .dinb(new_new_n1825__), .dout(new_new_n1005__));
  or1   g0474(.dina(new_new_n1888__), .dinb(new_new_n1830__), .dout(new_new_n1006__));
  or1   g0475(.dina(new_new_n1006__), .dinb(new_new_n558__), .dout(new_new_n1007__));
  or1   g0476(.dina(new_new_n1005__), .dinb(new_new_n559__), .dout(new_new_n1008__));
  and1  g0477(.dina(new_new_n1008__), .dinb(new_new_n1007__), .dout(new_new_n1009__));
  and1  g0478(.dina(new_new_n1886__), .dinb(new_new_n1835__), .dout(new_new_n1010__));
  or1   g0479(.dina(new_new_n1889__), .dinb(new_new_n1840__), .dout(new_new_n1011__));
  or1   g0480(.dina(new_new_n1011__), .dinb(new_new_n560__), .dout(new_new_n1012__));
  or1   g0481(.dina(new_new_n1010__), .dinb(new_new_n561__), .dout(new_new_n1013__));
  and1  g0482(.dina(new_new_n1013__), .dinb(new_new_n1012__), .dout(new_new_n1014__));
  and1  g0483(.dina(new_new_n1886__), .dinb(new_new_n1845__), .dout(new_new_n1015__));
  or1   g0484(.dina(new_new_n1889__), .dinb(new_new_n1850__), .dout(new_new_n1016__));
  or1   g0485(.dina(new_new_n1016__), .dinb(new_new_n562__), .dout(new_new_n1017__));
  or1   g0486(.dina(new_new_n1015__), .dinb(new_new_n563__), .dout(new_new_n1018__));
  and1  g0487(.dina(new_new_n1018__), .dinb(new_new_n1017__), .dout(new_new_n1019__));
  and1  g0488(.dina(new_new_n699__), .dinb(new_new_n1813__), .dout(new_new_n1020__));
  or1   g0489(.dina(new_new_n698__), .dinb(new_new_n1821__), .dout(new_new_n1021__));
  and1  g0490(.dina(new_new_n1020__), .dinb(new_new_n1836__), .dout(new_new_n1022__));
  or1   g0491(.dina(new_new_n1021__), .dinb(new_new_n1841__), .dout(new_new_n1023__));
  and1  g0492(.dina(new_new_n1022__), .dinb(new_new_n707__), .dout(new_new_n1024__));
  or1   g0493(.dina(new_new_n1023__), .dinb(new_new_n706__), .dout(new_new_n1025__));
  and1  g0494(.dina(new_new_n1024__), .dinb(new_new_n1891__), .dout(new_new_n1026__));
  or1   g0495(.dina(new_new_n1025__), .dinb(new_new_n1894__), .dout(new_new_n1027__));
  and1  g0496(.dina(new_new_n1897__), .dinb(new_new_n1783__), .dout(new_new_n1028__));
  or1   g0497(.dina(new_new_n1900__), .dinb(new_new_n1788__), .dout(new_new_n1029__));
  or1   g0498(.dina(new_new_n1029__), .dinb(new_new_n564__), .dout(new_new_n1030__));
  or1   g0499(.dina(new_new_n1028__), .dinb(new_new_n565__), .dout(new_new_n1031__));
  and1  g0500(.dina(new_new_n1031__), .dinb(new_new_n1030__), .dout(new_new_n1032__));
  and1  g0501(.dina(new_new_n1897__), .dinb(new_new_n1871__), .dout(new_new_n1033__));
  or1   g0502(.dina(new_new_n1900__), .dinb(new_new_n1876__), .dout(new_new_n1034__));
  or1   g0503(.dina(new_new_n1034__), .dinb(new_new_n566__), .dout(new_new_n1035__));
  or1   g0504(.dina(new_new_n1033__), .dinb(new_new_n567__), .dout(new_new_n1036__));
  and1  g0505(.dina(new_new_n1036__), .dinb(new_new_n1035__), .dout(new_new_n1037__));
  and1  g0506(.dina(new_new_n1898__), .dinb(new_new_n1793__), .dout(new_new_n1038__));
  or1   g0507(.dina(new_new_n1901__), .dinb(new_new_n1798__), .dout(new_new_n1039__));
  or1   g0508(.dina(new_new_n1039__), .dinb(new_new_n568__), .dout(new_new_n1040__));
  or1   g0509(.dina(new_new_n1038__), .dinb(new_new_n569__), .dout(new_new_n1041__));
  and1  g0510(.dina(new_new_n1041__), .dinb(new_new_n1040__), .dout(new_new_n1042__));
  and1  g0511(.dina(new_new_n1898__), .dinb(new_new_n1855__), .dout(new_new_n1043__));
  or1   g0512(.dina(new_new_n1901__), .dinb(new_new_n1860__), .dout(new_new_n1044__));
  or1   g0513(.dina(new_new_n1044__), .dinb(new_new_n570__), .dout(new_new_n1045__));
  or1   g0514(.dina(new_new_n1043__), .dinb(new_new_n571__), .dout(new_new_n1046__));
  and1  g0515(.dina(new_new_n1046__), .dinb(new_new_n1045__), .dout(new_new_n1047__));
  and1  g0516(.dina(new_new_n701__), .dinb(new_new_n1813__), .dout(new_new_n1048__));
  or1   g0517(.dina(new_new_n700__), .dinb(new_new_n1821__), .dout(new_new_n1049__));
  and1  g0518(.dina(new_new_n1048__), .dinb(new_new_n703__), .dout(new_new_n1050__));
  or1   g0519(.dina(new_new_n1049__), .dinb(new_new_n702__), .dout(new_new_n1051__));
  and1  g0520(.dina(new_new_n1050__), .dinb(new_new_n1846__), .dout(new_new_n1052__));
  or1   g0521(.dina(new_new_n1051__), .dinb(new_new_n1851__), .dout(new_new_n1053__));
  and1  g0522(.dina(new_new_n1052__), .dinb(new_new_n1891__), .dout(new_new_n1054__));
  or1   g0523(.dina(new_new_n1053__), .dinb(new_new_n1894__), .dout(new_new_n1055__));
  and1  g0524(.dina(new_new_n1903__), .dinb(new_new_n1783__), .dout(new_new_n1056__));
  or1   g0525(.dina(new_new_n1906__), .dinb(new_new_n1788__), .dout(new_new_n1057__));
  or1   g0526(.dina(new_new_n1057__), .dinb(new_new_n572__), .dout(new_new_n1058__));
  or1   g0527(.dina(new_new_n1056__), .dinb(new_new_n573__), .dout(new_new_n1059__));
  and1  g0528(.dina(new_new_n1059__), .dinb(new_new_n1058__), .dout(new_new_n1060__));
  and1  g0529(.dina(new_new_n1903__), .dinb(new_new_n1871__), .dout(new_new_n1061__));
  or1   g0530(.dina(new_new_n1906__), .dinb(new_new_n1876__), .dout(new_new_n1062__));
  or1   g0531(.dina(new_new_n1062__), .dinb(new_new_n574__), .dout(new_new_n1063__));
  or1   g0532(.dina(new_new_n1061__), .dinb(new_new_n575__), .dout(new_new_n1064__));
  and1  g0533(.dina(new_new_n1064__), .dinb(new_new_n1063__), .dout(new_new_n1065__));
  and1  g0534(.dina(new_new_n1904__), .dinb(new_new_n1793__), .dout(new_new_n1066__));
  or1   g0535(.dina(new_new_n1907__), .dinb(new_new_n1798__), .dout(new_new_n1067__));
  or1   g0536(.dina(new_new_n1067__), .dinb(new_new_n576__), .dout(new_new_n1068__));
  or1   g0537(.dina(new_new_n1066__), .dinb(new_new_n577__), .dout(new_new_n1069__));
  and1  g0538(.dina(new_new_n1069__), .dinb(new_new_n1068__), .dout(new_new_n1070__));
  and1  g0539(.dina(new_new_n1904__), .dinb(new_new_n1855__), .dout(new_new_n1071__));
  or1   g0540(.dina(new_new_n1907__), .dinb(new_new_n1860__), .dout(new_new_n1072__));
  or1   g0541(.dina(new_new_n1072__), .dinb(new_new_n578__), .dout(new_new_n1073__));
  or1   g0542(.dina(new_new_n1071__), .dinb(new_new_n579__), .dout(new_new_n1074__));
  and1  g0543(.dina(new_new_n1074__), .dinb(new_new_n1073__), .dout(new_new_n1075__));
  and1  g0544(.dina(new_new_n695__), .dinb(new_new_n1826__), .dout(new_new_n1076__));
  or1   g0545(.dina(new_new_n694__), .dinb(new_new_n1831__), .dout(new_new_n1077__));
  and1  g0546(.dina(new_new_n1076__), .dinb(new_new_n1836__), .dout(new_new_n1078__));
  or1   g0547(.dina(new_new_n1077__), .dinb(new_new_n1841__), .dout(new_new_n1079__));
  and1  g0548(.dina(new_new_n1078__), .dinb(new_new_n709__), .dout(new_new_n1080__));
  or1   g0549(.dina(new_new_n1079__), .dinb(new_new_n708__), .dout(new_new_n1081__));
  and1  g0550(.dina(new_new_n1080__), .dinb(new_new_n1892__), .dout(new_new_n1082__));
  or1   g0551(.dina(new_new_n1081__), .dinb(new_new_n1895__), .dout(new_new_n1083__));
  and1  g0552(.dina(new_new_n1909__), .dinb(new_new_n1784__), .dout(new_new_n1084__));
  or1   g0553(.dina(new_new_n1912__), .dinb(new_new_n1789__), .dout(new_new_n1085__));
  or1   g0554(.dina(new_new_n1085__), .dinb(new_new_n580__), .dout(new_new_n1086__));
  or1   g0555(.dina(new_new_n1084__), .dinb(new_new_n581__), .dout(new_new_n1087__));
  and1  g0556(.dina(new_new_n1087__), .dinb(new_new_n1086__), .dout(new_new_n1088__));
  and1  g0557(.dina(new_new_n1909__), .dinb(new_new_n1872__), .dout(new_new_n1089__));
  or1   g0558(.dina(new_new_n1912__), .dinb(new_new_n1877__), .dout(new_new_n1090__));
  or1   g0559(.dina(new_new_n1090__), .dinb(new_new_n582__), .dout(new_new_n1091__));
  or1   g0560(.dina(new_new_n1089__), .dinb(new_new_n583__), .dout(new_new_n1092__));
  and1  g0561(.dina(new_new_n1092__), .dinb(new_new_n1091__), .dout(new_new_n1093__));
  and1  g0562(.dina(new_new_n1910__), .dinb(new_new_n1794__), .dout(new_new_n1094__));
  or1   g0563(.dina(new_new_n1913__), .dinb(new_new_n1799__), .dout(new_new_n1095__));
  or1   g0564(.dina(new_new_n1095__), .dinb(new_new_n584__), .dout(new_new_n1096__));
  or1   g0565(.dina(new_new_n1094__), .dinb(new_new_n585__), .dout(new_new_n1097__));
  and1  g0566(.dina(new_new_n1097__), .dinb(new_new_n1096__), .dout(new_new_n1098__));
  and1  g0567(.dina(new_new_n1910__), .dinb(new_new_n1856__), .dout(new_new_n1099__));
  or1   g0568(.dina(new_new_n1913__), .dinb(new_new_n1861__), .dout(new_new_n1100__));
  or1   g0569(.dina(new_new_n1100__), .dinb(new_new_n586__), .dout(new_new_n1101__));
  or1   g0570(.dina(new_new_n1099__), .dinb(new_new_n587__), .dout(new_new_n1102__));
  and1  g0571(.dina(new_new_n1102__), .dinb(new_new_n1101__), .dout(new_new_n1103__));
  and1  g0572(.dina(new_new_n697__), .dinb(new_new_n1826__), .dout(new_new_n1104__));
  or1   g0573(.dina(new_new_n696__), .dinb(new_new_n1831__), .dout(new_new_n1105__));
  and1  g0574(.dina(new_new_n1104__), .dinb(new_new_n705__), .dout(new_new_n1106__));
  or1   g0575(.dina(new_new_n1105__), .dinb(new_new_n704__), .dout(new_new_n1107__));
  and1  g0576(.dina(new_new_n1106__), .dinb(new_new_n1846__), .dout(new_new_n1108__));
  or1   g0577(.dina(new_new_n1107__), .dinb(new_new_n1851__), .dout(new_new_n1109__));
  and1  g0578(.dina(new_new_n1108__), .dinb(new_new_n1892__), .dout(new_new_n1110__));
  or1   g0579(.dina(new_new_n1109__), .dinb(new_new_n1895__), .dout(new_new_n1111__));
  and1  g0580(.dina(new_new_n1915__), .dinb(new_new_n1784__), .dout(new_new_n1112__));
  or1   g0581(.dina(new_new_n1918__), .dinb(new_new_n1789__), .dout(new_new_n1113__));
  or1   g0582(.dina(new_new_n1113__), .dinb(new_new_n588__), .dout(new_new_n1114__));
  or1   g0583(.dina(new_new_n1112__), .dinb(new_new_n589__), .dout(new_new_n1115__));
  and1  g0584(.dina(new_new_n1115__), .dinb(new_new_n1114__), .dout(new_new_n1116__));
  and1  g0585(.dina(new_new_n1915__), .dinb(new_new_n1872__), .dout(new_new_n1117__));
  or1   g0586(.dina(new_new_n1918__), .dinb(new_new_n1877__), .dout(new_new_n1118__));
  or1   g0587(.dina(new_new_n1118__), .dinb(new_new_n590__), .dout(new_new_n1119__));
  or1   g0588(.dina(new_new_n1117__), .dinb(new_new_n591__), .dout(new_new_n1120__));
  and1  g0589(.dina(new_new_n1120__), .dinb(new_new_n1119__), .dout(new_new_n1121__));
  and1  g0590(.dina(new_new_n1916__), .dinb(new_new_n1794__), .dout(new_new_n1122__));
  or1   g0591(.dina(new_new_n1919__), .dinb(new_new_n1799__), .dout(new_new_n1123__));
  or1   g0592(.dina(new_new_n1123__), .dinb(new_new_n592__), .dout(new_new_n1124__));
  or1   g0593(.dina(new_new_n1122__), .dinb(new_new_n593__), .dout(new_new_n1125__));
  and1  g0594(.dina(new_new_n1125__), .dinb(new_new_n1124__), .dout(new_new_n1126__));
  and1  g0595(.dina(new_new_n1916__), .dinb(new_new_n1856__), .dout(new_new_n1127__));
  or1   g0596(.dina(new_new_n1919__), .dinb(new_new_n1861__), .dout(new_new_n1128__));
  or1   g0597(.dina(new_new_n1128__), .dinb(new_new_n594__), .dout(new_new_n1129__));
  or1   g0598(.dina(new_new_n1127__), .dinb(new_new_n595__), .dout(new_new_n1130__));
  and1  g0599(.dina(new_new_n1130__), .dinb(new_new_n1129__), .dout(new_new_n1131__));
  or1   g0600(.dina(new_new_n1920__), .dinb(new_new_n1921__), .dout(new_new_n1132__));
  or1   g0601(.dina(new_new_n1922__), .dinb(new_new_n1924__), .dout(new_new_n1133__));
  or1   g0602(.dina(new_new_n1133__), .dinb(new_new_n1926__), .dout(new_new_n1134__));
  or1   g0603(.dina(new_new_n1922__), .dinb(new_new_n1929__), .dout(new_new_n1135__));
  or1   g0604(.dina(new_new_n1135__), .dinb(new_new_n1932__), .dout(new_new_n1136__));
  or1   g0605(.dina(new_new_n1934__), .dinb(new_new_n1921__), .dout(new_new_n1137__));
  or1   g0606(.dina(new_new_n1137__), .dinb(new_new_n1924__), .dout(new_new_n1138__));
  or1   g0607(.dina(new_new_n1138__), .dinb(new_new_n1932__), .dout(new_new_n1139__));
  or1   g0608(.dina(new_new_n1920__), .dinb(new_new_n1937__), .dout(new_new_n1140__));
  or1   g0609(.dina(new_new_n1140__), .dinb(new_new_n1923__), .dout(new_new_n1141__));
  or1   g0610(.dina(new_new_n1141__), .dinb(new_new_n1931__), .dout(new_new_n1142__));
  and1  g0611(.dina(new_new_n1136__), .dinb(new_new_n1134__), .dout(new_new_n1143__));
  and1  g0612(.dina(new_new_n1143__), .dinb(new_new_n1139__), .dout(new_new_n1144__));
  and1  g0613(.dina(new_new_n1144__), .dinb(new_new_n1142__), .dout(new_new_n1145__));
  or1   g0614(.dina(new_new_n1939__), .dinb(new_new_n1940__), .dout(new_new_n1146__));
  or1   g0615(.dina(new_new_n1941__), .dinb(new_new_n1943__), .dout(new_new_n1147__));
  or1   g0616(.dina(new_new_n1147__), .dinb(new_new_n1945__), .dout(new_new_n1148__));
  or1   g0617(.dina(new_new_n1941__), .dinb(new_new_n1948__), .dout(new_new_n1149__));
  or1   g0618(.dina(new_new_n1149__), .dinb(new_new_n1951__), .dout(new_new_n1150__));
  or1   g0619(.dina(new_new_n1953__), .dinb(new_new_n1940__), .dout(new_new_n1151__));
  or1   g0620(.dina(new_new_n1151__), .dinb(new_new_n1943__), .dout(new_new_n1152__));
  or1   g0621(.dina(new_new_n1152__), .dinb(new_new_n1951__), .dout(new_new_n1153__));
  or1   g0622(.dina(new_new_n1939__), .dinb(new_new_n1956__), .dout(new_new_n1154__));
  or1   g0623(.dina(new_new_n1154__), .dinb(new_new_n1942__), .dout(new_new_n1155__));
  or1   g0624(.dina(new_new_n1155__), .dinb(new_new_n1950__), .dout(new_new_n1156__));
  and1  g0625(.dina(new_new_n1150__), .dinb(new_new_n1148__), .dout(new_new_n1157__));
  and1  g0626(.dina(new_new_n1157__), .dinb(new_new_n1153__), .dout(new_new_n1158__));
  and1  g0627(.dina(new_new_n1158__), .dinb(new_new_n1156__), .dout(new_new_n1159__));
  and1  g0628(.dina(new_new_n1958__), .dinb(new_new_n1960__), .dout(new_new_n1160__));
  or1   g0629(.dina(new_new_n1962__), .dinb(new_new_n1963__), .dout(new_new_n1161__));
  and1  g0630(.dina(new_new_n1962__), .dinb(new_new_n1963__), .dout(new_new_n1162__));
  or1   g0631(.dina(new_new_n1958__), .dinb(new_new_n1960__), .dout(new_new_n1163__));
  and1  g0632(.dina(new_new_n1163__), .dinb(new_new_n1161__), .dout(new_new_n1164__));
  or1   g0633(.dina(new_new_n1162__), .dinb(new_new_n1160__), .dout(new_new_n1165__));
  and1  g0634(.dina(new_new_n1964__), .dinb(new_new_n1966__), .dout(new_new_n1166__));
  or1   g0635(.dina(new_new_n1968__), .dinb(new_new_n1969__), .dout(new_new_n1167__));
  and1  g0636(.dina(new_new_n1968__), .dinb(new_new_n1969__), .dout(new_new_n1168__));
  or1   g0637(.dina(new_new_n1964__), .dinb(new_new_n1966__), .dout(new_new_n1169__));
  and1  g0638(.dina(new_new_n1169__), .dinb(new_new_n1167__), .dout(new_new_n1170__));
  or1   g0639(.dina(new_new_n1168__), .dinb(new_new_n1166__), .dout(new_new_n1171__));
  and1  g0640(.dina(new_new_n1970__), .dinb(new_new_n1971__), .dout(new_new_n1172__));
  or1   g0641(.dina(new_new_n1972__), .dinb(new_new_n1973__), .dout(new_new_n1173__));
  and1  g0642(.dina(new_new_n1972__), .dinb(new_new_n1973__), .dout(new_new_n1174__));
  or1   g0643(.dina(new_new_n1970__), .dinb(new_new_n1971__), .dout(new_new_n1175__));
  and1  g0644(.dina(new_new_n1175__), .dinb(new_new_n1173__), .dout(new_new_n1176__));
  or1   g0645(.dina(new_new_n1174__), .dinb(new_new_n1172__), .dout(new_new_n1177__));
  and1  g0646(.dina(new_new_n1976__), .dinb(new_new_n810__), .dout(new_new_n1178__));
  or1   g0647(.dina(new_new_n1983__), .dinb(new_new_n811__), .dout(new_new_n1179__));
  and1  g0648(.dina(new_new_n1989__), .dinb(new_new_n1992__), .dout(new_new_n1180__));
  or1   g0649(.dina(new_new_n1995__), .dinb(new_new_n1998__), .dout(new_new_n1181__));
  and1  g0650(.dina(new_new_n1995__), .dinb(new_new_n1998__), .dout(new_new_n1182__));
  or1   g0651(.dina(new_new_n1989__), .dinb(new_new_n1992__), .dout(new_new_n1183__));
  and1  g0652(.dina(new_new_n1183__), .dinb(new_new_n1181__), .dout(new_new_n1184__));
  or1   g0653(.dina(new_new_n1182__), .dinb(new_new_n1180__), .dout(new_new_n1185__));
  and1  g0654(.dina(new_new_n2000__), .dinb(new_new_n2001__), .dout(new_new_n1186__));
  or1   g0655(.dina(new_new_n2002__), .dinb(new_new_n2003__), .dout(new_new_n1187__));
  and1  g0656(.dina(new_new_n2002__), .dinb(new_new_n2003__), .dout(new_new_n1188__));
  or1   g0657(.dina(new_new_n2000__), .dinb(new_new_n2001__), .dout(new_new_n1189__));
  and1  g0658(.dina(new_new_n1189__), .dinb(new_new_n1187__), .dout(new_new_n1190__));
  or1   g0659(.dina(new_new_n1188__), .dinb(new_new_n1186__), .dout(new_new_n1191__));
  or1   g0660(.dina(new_new_n1190__), .dinb(new_new_n1177__), .dout(new_new_n1192__));
  or1   g0661(.dina(new_new_n1191__), .dinb(new_new_n1176__), .dout(new_new_n1193__));
  and1  g0662(.dina(new_new_n1193__), .dinb(new_new_n1192__), .dout(new_new_n1194__));
  and1  g0663(.dina(new_new_n2004__), .dinb(new_new_n2006__), .dout(new_new_n1195__));
  or1   g0664(.dina(new_new_n2008__), .dinb(new_new_n2009__), .dout(new_new_n1196__));
  and1  g0665(.dina(new_new_n2008__), .dinb(new_new_n2009__), .dout(new_new_n1197__));
  or1   g0666(.dina(new_new_n2004__), .dinb(new_new_n2006__), .dout(new_new_n1198__));
  and1  g0667(.dina(new_new_n1198__), .dinb(new_new_n1196__), .dout(new_new_n1199__));
  or1   g0668(.dina(new_new_n1197__), .dinb(new_new_n1195__), .dout(new_new_n1200__));
  and1  g0669(.dina(new_new_n2010__), .dinb(new_new_n2012__), .dout(new_new_n1201__));
  or1   g0670(.dina(new_new_n2014__), .dinb(new_new_n2015__), .dout(new_new_n1202__));
  and1  g0671(.dina(new_new_n2014__), .dinb(new_new_n2015__), .dout(new_new_n1203__));
  or1   g0672(.dina(new_new_n2010__), .dinb(new_new_n2012__), .dout(new_new_n1204__));
  and1  g0673(.dina(new_new_n1204__), .dinb(new_new_n1202__), .dout(new_new_n1205__));
  or1   g0674(.dina(new_new_n1203__), .dinb(new_new_n1201__), .dout(new_new_n1206__));
  and1  g0675(.dina(new_new_n2016__), .dinb(new_new_n2017__), .dout(new_new_n1207__));
  or1   g0676(.dina(new_new_n2018__), .dinb(new_new_n2019__), .dout(new_new_n1208__));
  and1  g0677(.dina(new_new_n2018__), .dinb(new_new_n2019__), .dout(new_new_n1209__));
  or1   g0678(.dina(new_new_n2016__), .dinb(new_new_n2017__), .dout(new_new_n1210__));
  and1  g0679(.dina(new_new_n1210__), .dinb(new_new_n1208__), .dout(new_new_n1211__));
  or1   g0680(.dina(new_new_n1209__), .dinb(new_new_n1207__), .dout(new_new_n1212__));
  and1  g0681(.dina(new_new_n1976__), .dinb(new_new_n812__), .dout(new_new_n1213__));
  or1   g0682(.dina(new_new_n1983__), .dinb(new_new_n813__), .dout(new_new_n1214__));
  and1  g0683(.dina(new_new_n2021__), .dinb(new_new_n2024__), .dout(new_new_n1215__));
  or1   g0684(.dina(new_new_n2027__), .dinb(new_new_n2030__), .dout(new_new_n1216__));
  and1  g0685(.dina(new_new_n2027__), .dinb(new_new_n2030__), .dout(new_new_n1217__));
  or1   g0686(.dina(new_new_n2021__), .dinb(new_new_n2024__), .dout(new_new_n1218__));
  and1  g0687(.dina(new_new_n1218__), .dinb(new_new_n1216__), .dout(new_new_n1219__));
  or1   g0688(.dina(new_new_n1217__), .dinb(new_new_n1215__), .dout(new_new_n1220__));
  and1  g0689(.dina(new_new_n2032__), .dinb(new_new_n2033__), .dout(new_new_n1221__));
  or1   g0690(.dina(new_new_n2034__), .dinb(new_new_n2035__), .dout(new_new_n1222__));
  and1  g0691(.dina(new_new_n2034__), .dinb(new_new_n2035__), .dout(new_new_n1223__));
  or1   g0692(.dina(new_new_n2032__), .dinb(new_new_n2033__), .dout(new_new_n1224__));
  and1  g0693(.dina(new_new_n1224__), .dinb(new_new_n1222__), .dout(new_new_n1225__));
  or1   g0694(.dina(new_new_n1223__), .dinb(new_new_n1221__), .dout(new_new_n1226__));
  or1   g0695(.dina(new_new_n1225__), .dinb(new_new_n1212__), .dout(new_new_n1227__));
  or1   g0696(.dina(new_new_n1226__), .dinb(new_new_n1211__), .dout(new_new_n1228__));
  and1  g0697(.dina(new_new_n1228__), .dinb(new_new_n1227__), .dout(new_new_n1229__));
  and1  g0698(.dina(new_new_n2036__), .dinb(new_new_n2038__), .dout(new_new_n1230__));
  or1   g0699(.dina(new_new_n2040__), .dinb(new_new_n2041__), .dout(new_new_n1231__));
  and1  g0700(.dina(new_new_n2040__), .dinb(new_new_n2041__), .dout(new_new_n1232__));
  or1   g0701(.dina(new_new_n2036__), .dinb(new_new_n2038__), .dout(new_new_n1233__));
  and1  g0702(.dina(new_new_n1233__), .dinb(new_new_n1231__), .dout(new_new_n1234__));
  or1   g0703(.dina(new_new_n1232__), .dinb(new_new_n1230__), .dout(new_new_n1235__));
  and1  g0704(.dina(new_new_n2042__), .dinb(new_new_n2044__), .dout(new_new_n1236__));
  or1   g0705(.dina(new_new_n2046__), .dinb(new_new_n2047__), .dout(new_new_n1237__));
  and1  g0706(.dina(new_new_n2046__), .dinb(new_new_n2047__), .dout(new_new_n1238__));
  or1   g0707(.dina(new_new_n2042__), .dinb(new_new_n2044__), .dout(new_new_n1239__));
  and1  g0708(.dina(new_new_n1239__), .dinb(new_new_n1237__), .dout(new_new_n1240__));
  or1   g0709(.dina(new_new_n1238__), .dinb(new_new_n1236__), .dout(new_new_n1241__));
  and1  g0710(.dina(new_new_n2048__), .dinb(new_new_n2049__), .dout(new_new_n1242__));
  or1   g0711(.dina(new_new_n2050__), .dinb(new_new_n2051__), .dout(new_new_n1243__));
  and1  g0712(.dina(new_new_n2050__), .dinb(new_new_n2051__), .dout(new_new_n1244__));
  or1   g0713(.dina(new_new_n2048__), .dinb(new_new_n2049__), .dout(new_new_n1245__));
  and1  g0714(.dina(new_new_n1245__), .dinb(new_new_n1243__), .dout(new_new_n1246__));
  or1   g0715(.dina(new_new_n1244__), .dinb(new_new_n1242__), .dout(new_new_n1247__));
  and1  g0716(.dina(new_new_n1977__), .dinb(new_new_n814__), .dout(new_new_n1248__));
  or1   g0717(.dina(new_new_n1984__), .dinb(new_new_n815__), .dout(new_new_n1249__));
  and1  g0718(.dina(new_new_n2031__), .dinb(new_new_n1993__), .dout(new_new_n1250__));
  or1   g0719(.dina(new_new_n2025__), .dinb(new_new_n1999__), .dout(new_new_n1251__));
  and1  g0720(.dina(new_new_n2025__), .dinb(new_new_n1999__), .dout(new_new_n1252__));
  or1   g0721(.dina(new_new_n2031__), .dinb(new_new_n1993__), .dout(new_new_n1253__));
  and1  g0722(.dina(new_new_n1253__), .dinb(new_new_n1251__), .dout(new_new_n1254__));
  or1   g0723(.dina(new_new_n1252__), .dinb(new_new_n1250__), .dout(new_new_n1255__));
  and1  g0724(.dina(new_new_n2052__), .dinb(new_new_n2053__), .dout(new_new_n1256__));
  or1   g0725(.dina(new_new_n2054__), .dinb(new_new_n2055__), .dout(new_new_n1257__));
  and1  g0726(.dina(new_new_n2054__), .dinb(new_new_n2055__), .dout(new_new_n1258__));
  or1   g0727(.dina(new_new_n2052__), .dinb(new_new_n2053__), .dout(new_new_n1259__));
  and1  g0728(.dina(new_new_n1259__), .dinb(new_new_n1257__), .dout(new_new_n1260__));
  or1   g0729(.dina(new_new_n1258__), .dinb(new_new_n1256__), .dout(new_new_n1261__));
  or1   g0730(.dina(new_new_n1260__), .dinb(new_new_n1247__), .dout(new_new_n1262__));
  or1   g0731(.dina(new_new_n1261__), .dinb(new_new_n1246__), .dout(new_new_n1263__));
  and1  g0732(.dina(new_new_n1263__), .dinb(new_new_n1262__), .dout(new_new_n1264__));
  and1  g0733(.dina(new_new_n2056__), .dinb(new_new_n2058__), .dout(new_new_n1265__));
  or1   g0734(.dina(new_new_n2060__), .dinb(new_new_n2061__), .dout(new_new_n1266__));
  and1  g0735(.dina(new_new_n2060__), .dinb(new_new_n2061__), .dout(new_new_n1267__));
  or1   g0736(.dina(new_new_n2056__), .dinb(new_new_n2058__), .dout(new_new_n1268__));
  and1  g0737(.dina(new_new_n1268__), .dinb(new_new_n1266__), .dout(new_new_n1269__));
  or1   g0738(.dina(new_new_n1267__), .dinb(new_new_n1265__), .dout(new_new_n1270__));
  and1  g0739(.dina(new_new_n2062__), .dinb(new_new_n2064__), .dout(new_new_n1271__));
  or1   g0740(.dina(new_new_n2066__), .dinb(new_new_n2067__), .dout(new_new_n1272__));
  and1  g0741(.dina(new_new_n2066__), .dinb(new_new_n2067__), .dout(new_new_n1273__));
  or1   g0742(.dina(new_new_n2062__), .dinb(new_new_n2064__), .dout(new_new_n1274__));
  and1  g0743(.dina(new_new_n1274__), .dinb(new_new_n1272__), .dout(new_new_n1275__));
  or1   g0744(.dina(new_new_n1273__), .dinb(new_new_n1271__), .dout(new_new_n1276__));
  and1  g0745(.dina(new_new_n2068__), .dinb(new_new_n2069__), .dout(new_new_n1277__));
  or1   g0746(.dina(new_new_n2070__), .dinb(new_new_n2071__), .dout(new_new_n1278__));
  and1  g0747(.dina(new_new_n2070__), .dinb(new_new_n2071__), .dout(new_new_n1279__));
  or1   g0748(.dina(new_new_n2068__), .dinb(new_new_n2069__), .dout(new_new_n1280__));
  and1  g0749(.dina(new_new_n1280__), .dinb(new_new_n1278__), .dout(new_new_n1281__));
  or1   g0750(.dina(new_new_n1279__), .dinb(new_new_n1277__), .dout(new_new_n1282__));
  and1  g0751(.dina(new_new_n1977__), .dinb(new_new_n816__), .dout(new_new_n1283__));
  or1   g0752(.dina(new_new_n1984__), .dinb(new_new_n817__), .dout(new_new_n1284__));
  and1  g0753(.dina(new_new_n2022__), .dinb(new_new_n1996__), .dout(new_new_n1285__));
  or1   g0754(.dina(new_new_n2028__), .dinb(new_new_n1990__), .dout(new_new_n1286__));
  and1  g0755(.dina(new_new_n2028__), .dinb(new_new_n1990__), .dout(new_new_n1287__));
  or1   g0756(.dina(new_new_n2022__), .dinb(new_new_n1996__), .dout(new_new_n1288__));
  and1  g0757(.dina(new_new_n1288__), .dinb(new_new_n1286__), .dout(new_new_n1289__));
  or1   g0758(.dina(new_new_n1287__), .dinb(new_new_n1285__), .dout(new_new_n1290__));
  and1  g0759(.dina(new_new_n2072__), .dinb(new_new_n2073__), .dout(new_new_n1291__));
  or1   g0760(.dina(new_new_n2074__), .dinb(new_new_n2075__), .dout(new_new_n1292__));
  and1  g0761(.dina(new_new_n2074__), .dinb(new_new_n2075__), .dout(new_new_n1293__));
  or1   g0762(.dina(new_new_n2072__), .dinb(new_new_n2073__), .dout(new_new_n1294__));
  and1  g0763(.dina(new_new_n1294__), .dinb(new_new_n1292__), .dout(new_new_n1295__));
  or1   g0764(.dina(new_new_n1293__), .dinb(new_new_n1291__), .dout(new_new_n1296__));
  or1   g0765(.dina(new_new_n1295__), .dinb(new_new_n1282__), .dout(new_new_n1297__));
  or1   g0766(.dina(new_new_n1296__), .dinb(new_new_n1281__), .dout(new_new_n1298__));
  and1  g0767(.dina(new_new_n1298__), .dinb(new_new_n1297__), .dout(new_new_n1299__));
  and1  g0768(.dina(new_new_n2076__), .dinb(new_new_n2078__), .dout(new_new_n1300__));
  or1   g0769(.dina(new_new_n2080__), .dinb(new_new_n2081__), .dout(new_new_n1301__));
  and1  g0770(.dina(new_new_n2080__), .dinb(new_new_n2081__), .dout(new_new_n1302__));
  or1   g0771(.dina(new_new_n2076__), .dinb(new_new_n2078__), .dout(new_new_n1303__));
  and1  g0772(.dina(new_new_n1303__), .dinb(new_new_n1301__), .dout(new_new_n1304__));
  or1   g0773(.dina(new_new_n1302__), .dinb(new_new_n1300__), .dout(new_new_n1305__));
  and1  g0774(.dina(new_new_n2082__), .dinb(new_new_n2084__), .dout(new_new_n1306__));
  or1   g0775(.dina(new_new_n2086__), .dinb(new_new_n2087__), .dout(new_new_n1307__));
  and1  g0776(.dina(new_new_n2086__), .dinb(new_new_n2087__), .dout(new_new_n1308__));
  or1   g0777(.dina(new_new_n2082__), .dinb(new_new_n2084__), .dout(new_new_n1309__));
  and1  g0778(.dina(new_new_n1309__), .dinb(new_new_n1307__), .dout(new_new_n1310__));
  or1   g0779(.dina(new_new_n1308__), .dinb(new_new_n1306__), .dout(new_new_n1311__));
  and1  g0780(.dina(new_new_n2088__), .dinb(new_new_n2089__), .dout(new_new_n1312__));
  or1   g0781(.dina(new_new_n2090__), .dinb(new_new_n2091__), .dout(new_new_n1313__));
  and1  g0782(.dina(new_new_n2090__), .dinb(new_new_n2091__), .dout(new_new_n1314__));
  or1   g0783(.dina(new_new_n2088__), .dinb(new_new_n2089__), .dout(new_new_n1315__));
  and1  g0784(.dina(new_new_n1315__), .dinb(new_new_n1313__), .dout(new_new_n1316__));
  or1   g0785(.dina(new_new_n1314__), .dinb(new_new_n1312__), .dout(new_new_n1317__));
  and1  g0786(.dina(new_new_n1979__), .dinb(new_new_n818__), .dout(new_new_n1318__));
  or1   g0787(.dina(new_new_n1986__), .dinb(new_new_n819__), .dout(new_new_n1319__));
  and1  g0788(.dina(new_new_n2093__), .dinb(new_new_n2096__), .dout(new_new_n1320__));
  or1   g0789(.dina(new_new_n2099__), .dinb(new_new_n2102__), .dout(new_new_n1321__));
  and1  g0790(.dina(new_new_n2099__), .dinb(new_new_n2102__), .dout(new_new_n1322__));
  or1   g0791(.dina(new_new_n2093__), .dinb(new_new_n2096__), .dout(new_new_n1323__));
  and1  g0792(.dina(new_new_n1323__), .dinb(new_new_n1321__), .dout(new_new_n1324__));
  or1   g0793(.dina(new_new_n1322__), .dinb(new_new_n1320__), .dout(new_new_n1325__));
  and1  g0794(.dina(new_new_n2104__), .dinb(new_new_n2105__), .dout(new_new_n1326__));
  or1   g0795(.dina(new_new_n2106__), .dinb(new_new_n2107__), .dout(new_new_n1327__));
  and1  g0796(.dina(new_new_n2106__), .dinb(new_new_n2107__), .dout(new_new_n1328__));
  or1   g0797(.dina(new_new_n2104__), .dinb(new_new_n2105__), .dout(new_new_n1329__));
  and1  g0798(.dina(new_new_n1329__), .dinb(new_new_n1327__), .dout(new_new_n1330__));
  or1   g0799(.dina(new_new_n1328__), .dinb(new_new_n1326__), .dout(new_new_n1331__));
  or1   g0800(.dina(new_new_n1330__), .dinb(new_new_n1317__), .dout(new_new_n1332__));
  or1   g0801(.dina(new_new_n1331__), .dinb(new_new_n1316__), .dout(new_new_n1333__));
  and1  g0802(.dina(new_new_n1333__), .dinb(new_new_n1332__), .dout(new_new_n1334__));
  and1  g0803(.dina(new_new_n2108__), .dinb(new_new_n2110__), .dout(new_new_n1335__));
  or1   g0804(.dina(new_new_n2112__), .dinb(new_new_n2113__), .dout(new_new_n1336__));
  and1  g0805(.dina(new_new_n2112__), .dinb(new_new_n2113__), .dout(new_new_n1337__));
  or1   g0806(.dina(new_new_n2108__), .dinb(new_new_n2110__), .dout(new_new_n1338__));
  and1  g0807(.dina(new_new_n1338__), .dinb(new_new_n1336__), .dout(new_new_n1339__));
  or1   g0808(.dina(new_new_n1337__), .dinb(new_new_n1335__), .dout(new_new_n1340__));
  and1  g0809(.dina(new_new_n2114__), .dinb(new_new_n2116__), .dout(new_new_n1341__));
  or1   g0810(.dina(new_new_n2118__), .dinb(new_new_n2119__), .dout(new_new_n1342__));
  and1  g0811(.dina(new_new_n2118__), .dinb(new_new_n2119__), .dout(new_new_n1343__));
  or1   g0812(.dina(new_new_n2114__), .dinb(new_new_n2116__), .dout(new_new_n1344__));
  and1  g0813(.dina(new_new_n1344__), .dinb(new_new_n1342__), .dout(new_new_n1345__));
  or1   g0814(.dina(new_new_n1343__), .dinb(new_new_n1341__), .dout(new_new_n1346__));
  and1  g0815(.dina(new_new_n2120__), .dinb(new_new_n2121__), .dout(new_new_n1347__));
  or1   g0816(.dina(new_new_n2122__), .dinb(new_new_n2123__), .dout(new_new_n1348__));
  and1  g0817(.dina(new_new_n2122__), .dinb(new_new_n2123__), .dout(new_new_n1349__));
  or1   g0818(.dina(new_new_n2120__), .dinb(new_new_n2121__), .dout(new_new_n1350__));
  and1  g0819(.dina(new_new_n1350__), .dinb(new_new_n1348__), .dout(new_new_n1351__));
  or1   g0820(.dina(new_new_n1349__), .dinb(new_new_n1347__), .dout(new_new_n1352__));
  and1  g0821(.dina(new_new_n1979__), .dinb(new_new_n820__), .dout(new_new_n1353__));
  or1   g0822(.dina(new_new_n1986__), .dinb(new_new_n821__), .dout(new_new_n1354__));
  and1  g0823(.dina(new_new_n2125__), .dinb(new_new_n2128__), .dout(new_new_n1355__));
  or1   g0824(.dina(new_new_n2131__), .dinb(new_new_n2134__), .dout(new_new_n1356__));
  and1  g0825(.dina(new_new_n2131__), .dinb(new_new_n2134__), .dout(new_new_n1357__));
  or1   g0826(.dina(new_new_n2125__), .dinb(new_new_n2128__), .dout(new_new_n1358__));
  and1  g0827(.dina(new_new_n1358__), .dinb(new_new_n1356__), .dout(new_new_n1359__));
  or1   g0828(.dina(new_new_n1357__), .dinb(new_new_n1355__), .dout(new_new_n1360__));
  and1  g0829(.dina(new_new_n2136__), .dinb(new_new_n2137__), .dout(new_new_n1361__));
  or1   g0830(.dina(new_new_n2138__), .dinb(new_new_n2139__), .dout(new_new_n1362__));
  and1  g0831(.dina(new_new_n2138__), .dinb(new_new_n2139__), .dout(new_new_n1363__));
  or1   g0832(.dina(new_new_n2136__), .dinb(new_new_n2137__), .dout(new_new_n1364__));
  and1  g0833(.dina(new_new_n1364__), .dinb(new_new_n1362__), .dout(new_new_n1365__));
  or1   g0834(.dina(new_new_n1363__), .dinb(new_new_n1361__), .dout(new_new_n1366__));
  or1   g0835(.dina(new_new_n1365__), .dinb(new_new_n1352__), .dout(new_new_n1367__));
  or1   g0836(.dina(new_new_n1366__), .dinb(new_new_n1351__), .dout(new_new_n1368__));
  and1  g0837(.dina(new_new_n1368__), .dinb(new_new_n1367__), .dout(new_new_n1369__));
  and1  g0838(.dina(new_new_n2140__), .dinb(new_new_n2142__), .dout(new_new_n1370__));
  or1   g0839(.dina(new_new_n2144__), .dinb(new_new_n2145__), .dout(new_new_n1371__));
  and1  g0840(.dina(new_new_n2144__), .dinb(new_new_n2145__), .dout(new_new_n1372__));
  or1   g0841(.dina(new_new_n2140__), .dinb(new_new_n2142__), .dout(new_new_n1373__));
  and1  g0842(.dina(new_new_n1373__), .dinb(new_new_n1371__), .dout(new_new_n1374__));
  or1   g0843(.dina(new_new_n1372__), .dinb(new_new_n1370__), .dout(new_new_n1375__));
  and1  g0844(.dina(new_new_n2146__), .dinb(new_new_n2148__), .dout(new_new_n1376__));
  or1   g0845(.dina(new_new_n2150__), .dinb(new_new_n2151__), .dout(new_new_n1377__));
  and1  g0846(.dina(new_new_n2150__), .dinb(new_new_n2151__), .dout(new_new_n1378__));
  or1   g0847(.dina(new_new_n2146__), .dinb(new_new_n2148__), .dout(new_new_n1379__));
  and1  g0848(.dina(new_new_n1379__), .dinb(new_new_n1377__), .dout(new_new_n1380__));
  or1   g0849(.dina(new_new_n1378__), .dinb(new_new_n1376__), .dout(new_new_n1381__));
  and1  g0850(.dina(new_new_n2152__), .dinb(new_new_n2153__), .dout(new_new_n1382__));
  or1   g0851(.dina(new_new_n2154__), .dinb(new_new_n2155__), .dout(new_new_n1383__));
  and1  g0852(.dina(new_new_n2154__), .dinb(new_new_n2155__), .dout(new_new_n1384__));
  or1   g0853(.dina(new_new_n2152__), .dinb(new_new_n2153__), .dout(new_new_n1385__));
  and1  g0854(.dina(new_new_n1385__), .dinb(new_new_n1383__), .dout(new_new_n1386__));
  or1   g0855(.dina(new_new_n1384__), .dinb(new_new_n1382__), .dout(new_new_n1387__));
  and1  g0856(.dina(new_new_n1980__), .dinb(new_new_n822__), .dout(new_new_n1388__));
  or1   g0857(.dina(new_new_n1987__), .dinb(new_new_n823__), .dout(new_new_n1389__));
  and1  g0858(.dina(new_new_n2135__), .dinb(new_new_n2097__), .dout(new_new_n1390__));
  or1   g0859(.dina(new_new_n2129__), .dinb(new_new_n2103__), .dout(new_new_n1391__));
  and1  g0860(.dina(new_new_n2129__), .dinb(new_new_n2103__), .dout(new_new_n1392__));
  or1   g0861(.dina(new_new_n2135__), .dinb(new_new_n2097__), .dout(new_new_n1393__));
  and1  g0862(.dina(new_new_n1393__), .dinb(new_new_n1391__), .dout(new_new_n1394__));
  or1   g0863(.dina(new_new_n1392__), .dinb(new_new_n1390__), .dout(new_new_n1395__));
  and1  g0864(.dina(new_new_n2156__), .dinb(new_new_n2157__), .dout(new_new_n1396__));
  or1   g0865(.dina(new_new_n2158__), .dinb(new_new_n2159__), .dout(new_new_n1397__));
  and1  g0866(.dina(new_new_n2158__), .dinb(new_new_n2159__), .dout(new_new_n1398__));
  or1   g0867(.dina(new_new_n2156__), .dinb(new_new_n2157__), .dout(new_new_n1399__));
  and1  g0868(.dina(new_new_n1399__), .dinb(new_new_n1397__), .dout(new_new_n1400__));
  or1   g0869(.dina(new_new_n1398__), .dinb(new_new_n1396__), .dout(new_new_n1401__));
  or1   g0870(.dina(new_new_n1400__), .dinb(new_new_n1387__), .dout(new_new_n1402__));
  or1   g0871(.dina(new_new_n1401__), .dinb(new_new_n1386__), .dout(new_new_n1403__));
  and1  g0872(.dina(new_new_n1403__), .dinb(new_new_n1402__), .dout(new_new_n1404__));
  and1  g0873(.dina(new_new_n2160__), .dinb(new_new_n2162__), .dout(new_new_n1405__));
  or1   g0874(.dina(new_new_n2164__), .dinb(new_new_n2165__), .dout(new_new_n1406__));
  and1  g0875(.dina(new_new_n2164__), .dinb(new_new_n2165__), .dout(new_new_n1407__));
  or1   g0876(.dina(new_new_n2160__), .dinb(new_new_n2162__), .dout(new_new_n1408__));
  and1  g0877(.dina(new_new_n1408__), .dinb(new_new_n1406__), .dout(new_new_n1409__));
  or1   g0878(.dina(new_new_n1407__), .dinb(new_new_n1405__), .dout(new_new_n1410__));
  and1  g0879(.dina(new_new_n2166__), .dinb(new_new_n2168__), .dout(new_new_n1411__));
  or1   g0880(.dina(new_new_n2170__), .dinb(new_new_n2171__), .dout(new_new_n1412__));
  and1  g0881(.dina(new_new_n2170__), .dinb(new_new_n2171__), .dout(new_new_n1413__));
  or1   g0882(.dina(new_new_n2166__), .dinb(new_new_n2168__), .dout(new_new_n1414__));
  and1  g0883(.dina(new_new_n1414__), .dinb(new_new_n1412__), .dout(new_new_n1415__));
  or1   g0884(.dina(new_new_n1413__), .dinb(new_new_n1411__), .dout(new_new_n1416__));
  and1  g0885(.dina(new_new_n2172__), .dinb(new_new_n2173__), .dout(new_new_n1417__));
  or1   g0886(.dina(new_new_n2174__), .dinb(new_new_n2175__), .dout(new_new_n1418__));
  and1  g0887(.dina(new_new_n2174__), .dinb(new_new_n2175__), .dout(new_new_n1419__));
  or1   g0888(.dina(new_new_n2172__), .dinb(new_new_n2173__), .dout(new_new_n1420__));
  and1  g0889(.dina(new_new_n1420__), .dinb(new_new_n1418__), .dout(new_new_n1421__));
  or1   g0890(.dina(new_new_n1419__), .dinb(new_new_n1417__), .dout(new_new_n1422__));
  and1  g0891(.dina(new_new_n1980__), .dinb(new_new_n824__), .dout(new_new_n1423__));
  or1   g0892(.dina(new_new_n1987__), .dinb(new_new_n825__), .dout(new_new_n1424__));
  and1  g0893(.dina(new_new_n2126__), .dinb(new_new_n2100__), .dout(new_new_n1425__));
  or1   g0894(.dina(new_new_n2132__), .dinb(new_new_n2094__), .dout(new_new_n1426__));
  and1  g0895(.dina(new_new_n2132__), .dinb(new_new_n2094__), .dout(new_new_n1427__));
  or1   g0896(.dina(new_new_n2126__), .dinb(new_new_n2100__), .dout(new_new_n1428__));
  and1  g0897(.dina(new_new_n1428__), .dinb(new_new_n1426__), .dout(new_new_n1429__));
  or1   g0898(.dina(new_new_n1427__), .dinb(new_new_n1425__), .dout(new_new_n1430__));
  and1  g0899(.dina(new_new_n2176__), .dinb(new_new_n2177__), .dout(new_new_n1431__));
  or1   g0900(.dina(new_new_n2178__), .dinb(new_new_n2179__), .dout(new_new_n1432__));
  and1  g0901(.dina(new_new_n2178__), .dinb(new_new_n2179__), .dout(new_new_n1433__));
  or1   g0902(.dina(new_new_n2176__), .dinb(new_new_n2177__), .dout(new_new_n1434__));
  and1  g0903(.dina(new_new_n1434__), .dinb(new_new_n1432__), .dout(new_new_n1435__));
  or1   g0904(.dina(new_new_n1433__), .dinb(new_new_n1431__), .dout(new_new_n1436__));
  or1   g0905(.dina(new_new_n1435__), .dinb(new_new_n1422__), .dout(new_new_n1437__));
  or1   g0906(.dina(new_new_n1436__), .dinb(new_new_n1421__), .dout(new_new_n1438__));
  and1  g0907(.dina(new_new_n1438__), .dinb(new_new_n1437__), .dout(new_new_n1439__));
  and1  g0908(.dina(new_new_n2180__), .dinb(new_new_n2182__), .dout(new_new_n1440__));
  or1   g0909(.dina(new_new_n2184__), .dinb(new_new_n2185__), .dout(new_new_n1441__));
  and1  g0910(.dina(new_new_n2184__), .dinb(new_new_n2185__), .dout(new_new_n1442__));
  or1   g0911(.dina(new_new_n2180__), .dinb(new_new_n2182__), .dout(new_new_n1443__));
  and1  g0912(.dina(new_new_n1443__), .dinb(new_new_n1441__), .dout(new_new_n1444__));
  or1   g0913(.dina(new_new_n1442__), .dinb(new_new_n1440__), .dout(new_new_n1445__));
  and1  g0914(.dina(new_new_n2186__), .dinb(new_new_n2188__), .dout(new_new_n1446__));
  or1   g0915(.dina(new_new_n2190__), .dinb(new_new_n2191__), .dout(new_new_n1447__));
  and1  g0916(.dina(new_new_n2190__), .dinb(new_new_n2191__), .dout(new_new_n1448__));
  or1   g0917(.dina(new_new_n2186__), .dinb(new_new_n2188__), .dout(new_new_n1449__));
  and1  g0918(.dina(new_new_n1449__), .dinb(new_new_n1447__), .dout(new_new_n1450__));
  or1   g0919(.dina(new_new_n1448__), .dinb(new_new_n1446__), .dout(new_new_n1451__));
  or1   g0920(.dina(new_new_n1450__), .dinb(new_new_n1445__), .dout(new_new_n1452__));
  or1   g0921(.dina(new_new_n1451__), .dinb(new_new_n1444__), .dout(new_new_n1453__));
  and1  g0922(.dina(new_new_n1453__), .dinb(new_new_n1452__), .dout(new_new_n1454__));
  and1  g0923(.dina(new_new_n2192__), .dinb(new_new_n2194__), .dout(new_new_n1455__));
  or1   g0924(.dina(new_new_n2196__), .dinb(new_new_n2197__), .dout(new_new_n1456__));
  and1  g0925(.dina(new_new_n2196__), .dinb(new_new_n2197__), .dout(new_new_n1457__));
  or1   g0926(.dina(new_new_n2192__), .dinb(new_new_n2194__), .dout(new_new_n1458__));
  and1  g0927(.dina(new_new_n1458__), .dinb(new_new_n1456__), .dout(new_new_n1459__));
  or1   g0928(.dina(new_new_n1457__), .dinb(new_new_n1455__), .dout(new_new_n1460__));
  and1  g0929(.dina(new_new_n2198__), .dinb(new_new_n2200__), .dout(new_new_n1461__));
  or1   g0930(.dina(new_new_n2202__), .dinb(new_new_n2203__), .dout(new_new_n1462__));
  and1  g0931(.dina(new_new_n2202__), .dinb(new_new_n2203__), .dout(new_new_n1463__));
  or1   g0932(.dina(new_new_n2198__), .dinb(new_new_n2200__), .dout(new_new_n1464__));
  and1  g0933(.dina(new_new_n1464__), .dinb(new_new_n1462__), .dout(new_new_n1465__));
  or1   g0934(.dina(new_new_n1463__), .dinb(new_new_n1461__), .dout(new_new_n1466__));
  or1   g0935(.dina(new_new_n1465__), .dinb(new_new_n1460__), .dout(new_new_n1467__));
  or1   g0936(.dina(new_new_n1466__), .dinb(new_new_n1459__), .dout(new_new_n1468__));
  and1  g0937(.dina(new_new_n1468__), .dinb(new_new_n1467__), .dout(new_new_n1469__));
  and1  g0938(.dina(new_new_n2204__), .dinb(new_new_n2206__), .dout(new_new_n1470__));
  or1   g0939(.dina(new_new_n2208__), .dinb(new_new_n2209__), .dout(new_new_n1471__));
  and1  g0940(.dina(new_new_n2208__), .dinb(new_new_n2209__), .dout(new_new_n1472__));
  or1   g0941(.dina(new_new_n2204__), .dinb(new_new_n2206__), .dout(new_new_n1473__));
  and1  g0942(.dina(new_new_n1473__), .dinb(new_new_n1471__), .dout(new_new_n1474__));
  or1   g0943(.dina(new_new_n1472__), .dinb(new_new_n1470__), .dout(new_new_n1475__));
  and1  g0944(.dina(new_new_n2210__), .dinb(new_new_n2212__), .dout(new_new_n1476__));
  or1   g0945(.dina(new_new_n2214__), .dinb(new_new_n2215__), .dout(new_new_n1477__));
  and1  g0946(.dina(new_new_n2214__), .dinb(new_new_n2215__), .dout(new_new_n1478__));
  or1   g0947(.dina(new_new_n2210__), .dinb(new_new_n2212__), .dout(new_new_n1479__));
  and1  g0948(.dina(new_new_n1479__), .dinb(new_new_n1477__), .dout(new_new_n1480__));
  or1   g0949(.dina(new_new_n1478__), .dinb(new_new_n1476__), .dout(new_new_n1481__));
  or1   g0950(.dina(new_new_n1480__), .dinb(new_new_n1475__), .dout(new_new_n1482__));
  or1   g0951(.dina(new_new_n1481__), .dinb(new_new_n1474__), .dout(new_new_n1483__));
  and1  g0952(.dina(new_new_n1483__), .dinb(new_new_n1482__), .dout(new_new_n1484__));
  and1  g0953(.dina(new_new_n2216__), .dinb(new_new_n2218__), .dout(new_new_n1485__));
  or1   g0954(.dina(new_new_n2220__), .dinb(new_new_n2221__), .dout(new_new_n1486__));
  and1  g0955(.dina(new_new_n2220__), .dinb(new_new_n2221__), .dout(new_new_n1487__));
  or1   g0956(.dina(new_new_n2216__), .dinb(new_new_n2218__), .dout(new_new_n1488__));
  and1  g0957(.dina(new_new_n1488__), .dinb(new_new_n1486__), .dout(new_new_n1489__));
  or1   g0958(.dina(new_new_n1487__), .dinb(new_new_n1485__), .dout(new_new_n1490__));
  and1  g0959(.dina(new_new_n2222__), .dinb(new_new_n2224__), .dout(new_new_n1491__));
  or1   g0960(.dina(new_new_n2226__), .dinb(new_new_n2227__), .dout(new_new_n1492__));
  and1  g0961(.dina(new_new_n2226__), .dinb(new_new_n2227__), .dout(new_new_n1493__));
  or1   g0962(.dina(new_new_n2222__), .dinb(new_new_n2224__), .dout(new_new_n1494__));
  and1  g0963(.dina(new_new_n1494__), .dinb(new_new_n1492__), .dout(new_new_n1495__));
  or1   g0964(.dina(new_new_n1493__), .dinb(new_new_n1491__), .dout(new_new_n1496__));
  or1   g0965(.dina(new_new_n1495__), .dinb(new_new_n1490__), .dout(new_new_n1497__));
  or1   g0966(.dina(new_new_n1496__), .dinb(new_new_n1489__), .dout(new_new_n1498__));
  and1  g0967(.dina(new_new_n1498__), .dinb(new_new_n1497__), .dout(new_new_n1499__));
  and1  g0968(.dina(new_new_n2228__), .dinb(new_new_n2230__), .dout(new_new_n1500__));
  or1   g0969(.dina(new_new_n2232__), .dinb(new_new_n2233__), .dout(new_new_n1501__));
  and1  g0970(.dina(new_new_n2232__), .dinb(new_new_n2233__), .dout(new_new_n1502__));
  or1   g0971(.dina(new_new_n2228__), .dinb(new_new_n2230__), .dout(new_new_n1503__));
  and1  g0972(.dina(new_new_n1503__), .dinb(new_new_n1501__), .dout(new_new_n1504__));
  or1   g0973(.dina(new_new_n1502__), .dinb(new_new_n1500__), .dout(new_new_n1505__));
  and1  g0974(.dina(new_new_n2234__), .dinb(new_new_n2236__), .dout(new_new_n1506__));
  or1   g0975(.dina(new_new_n2238__), .dinb(new_new_n2239__), .dout(new_new_n1507__));
  and1  g0976(.dina(new_new_n2238__), .dinb(new_new_n2239__), .dout(new_new_n1508__));
  or1   g0977(.dina(new_new_n2234__), .dinb(new_new_n2236__), .dout(new_new_n1509__));
  and1  g0978(.dina(new_new_n1509__), .dinb(new_new_n1507__), .dout(new_new_n1510__));
  or1   g0979(.dina(new_new_n1508__), .dinb(new_new_n1506__), .dout(new_new_n1511__));
  or1   g0980(.dina(new_new_n1510__), .dinb(new_new_n1505__), .dout(new_new_n1512__));
  or1   g0981(.dina(new_new_n1511__), .dinb(new_new_n1504__), .dout(new_new_n1513__));
  and1  g0982(.dina(new_new_n1513__), .dinb(new_new_n1512__), .dout(new_new_n1514__));
  and1  g0983(.dina(new_new_n2240__), .dinb(new_new_n2242__), .dout(new_new_n1515__));
  or1   g0984(.dina(new_new_n2244__), .dinb(new_new_n2245__), .dout(new_new_n1516__));
  and1  g0985(.dina(new_new_n2244__), .dinb(new_new_n2245__), .dout(new_new_n1517__));
  or1   g0986(.dina(new_new_n2240__), .dinb(new_new_n2242__), .dout(new_new_n1518__));
  and1  g0987(.dina(new_new_n1518__), .dinb(new_new_n1516__), .dout(new_new_n1519__));
  or1   g0988(.dina(new_new_n1517__), .dinb(new_new_n1515__), .dout(new_new_n1520__));
  and1  g0989(.dina(new_new_n2246__), .dinb(new_new_n2248__), .dout(new_new_n1521__));
  or1   g0990(.dina(new_new_n2250__), .dinb(new_new_n2251__), .dout(new_new_n1522__));
  and1  g0991(.dina(new_new_n2250__), .dinb(new_new_n2251__), .dout(new_new_n1523__));
  or1   g0992(.dina(new_new_n2246__), .dinb(new_new_n2248__), .dout(new_new_n1524__));
  and1  g0993(.dina(new_new_n1524__), .dinb(new_new_n1522__), .dout(new_new_n1525__));
  or1   g0994(.dina(new_new_n1523__), .dinb(new_new_n1521__), .dout(new_new_n1526__));
  or1   g0995(.dina(new_new_n1525__), .dinb(new_new_n1520__), .dout(new_new_n1527__));
  or1   g0996(.dina(new_new_n1526__), .dinb(new_new_n1519__), .dout(new_new_n1528__));
  and1  g0997(.dina(new_new_n1528__), .dinb(new_new_n1527__), .dout(new_new_n1529__));
  and1  g0998(.dina(new_new_n2252__), .dinb(new_new_n2254__), .dout(new_new_n1530__));
  or1   g0999(.dina(new_new_n2256__), .dinb(new_new_n2257__), .dout(new_new_n1531__));
  and1  g1000(.dina(new_new_n2256__), .dinb(new_new_n2257__), .dout(new_new_n1532__));
  or1   g1001(.dina(new_new_n2252__), .dinb(new_new_n2254__), .dout(new_new_n1533__));
  and1  g1002(.dina(new_new_n1533__), .dinb(new_new_n1531__), .dout(new_new_n1534__));
  or1   g1003(.dina(new_new_n1532__), .dinb(new_new_n1530__), .dout(new_new_n1535__));
  and1  g1004(.dina(new_new_n2258__), .dinb(new_new_n2260__), .dout(new_new_n1536__));
  or1   g1005(.dina(new_new_n2262__), .dinb(new_new_n2263__), .dout(new_new_n1537__));
  and1  g1006(.dina(new_new_n2262__), .dinb(new_new_n2263__), .dout(new_new_n1538__));
  or1   g1007(.dina(new_new_n2258__), .dinb(new_new_n2260__), .dout(new_new_n1539__));
  and1  g1008(.dina(new_new_n1539__), .dinb(new_new_n1537__), .dout(new_new_n1540__));
  or1   g1009(.dina(new_new_n1538__), .dinb(new_new_n1536__), .dout(new_new_n1541__));
  or1   g1010(.dina(new_new_n1540__), .dinb(new_new_n1535__), .dout(new_new_n1542__));
  or1   g1011(.dina(new_new_n1541__), .dinb(new_new_n1534__), .dout(new_new_n1543__));
  and1  g1012(.dina(new_new_n1543__), .dinb(new_new_n1542__), .dout(new_new_n1544__));
  and1  g1013(.dina(new_new_n2264__), .dinb(new_new_n2266__), .dout(new_new_n1545__));
  or1   g1014(.dina(new_new_n2268__), .dinb(new_new_n2269__), .dout(new_new_n1546__));
  and1  g1015(.dina(new_new_n2268__), .dinb(new_new_n2269__), .dout(new_new_n1547__));
  or1   g1016(.dina(new_new_n2264__), .dinb(new_new_n2266__), .dout(new_new_n1548__));
  and1  g1017(.dina(new_new_n1548__), .dinb(new_new_n1546__), .dout(new_new_n1549__));
  or1   g1018(.dina(new_new_n1547__), .dinb(new_new_n1545__), .dout(new_new_n1550__));
  and1  g1019(.dina(new_new_n2270__), .dinb(new_new_n2272__), .dout(new_new_n1551__));
  or1   g1020(.dina(new_new_n2274__), .dinb(new_new_n2275__), .dout(new_new_n1552__));
  and1  g1021(.dina(new_new_n2274__), .dinb(new_new_n2275__), .dout(new_new_n1553__));
  or1   g1022(.dina(new_new_n2270__), .dinb(new_new_n2272__), .dout(new_new_n1554__));
  and1  g1023(.dina(new_new_n1554__), .dinb(new_new_n1552__), .dout(new_new_n1555__));
  or1   g1024(.dina(new_new_n1553__), .dinb(new_new_n1551__), .dout(new_new_n1556__));
  or1   g1025(.dina(new_new_n1555__), .dinb(new_new_n1550__), .dout(new_new_n1557__));
  or1   g1026(.dina(new_new_n1556__), .dinb(new_new_n1549__), .dout(new_new_n1558__));
  and1  g1027(.dina(new_new_n1558__), .dinb(new_new_n1557__), .dout(new_new_n1559__));
  not1  g1028(.din(new_new_n920__), .dout(G468));
  not1  g1029(.din(new_new_n925__), .dout(G469));
  not1  g1030(.din(new_new_n930__), .dout(G470));
  not1  g1031(.din(new_new_n935__), .dout(G471));
  not1  g1032(.din(new_new_n948__), .dout(G472));
  not1  g1033(.din(new_new_n953__), .dout(G473));
  not1  g1034(.din(new_new_n958__), .dout(G474));
  not1  g1035(.din(new_new_n963__), .dout(G475));
  not1  g1036(.din(new_new_n976__), .dout(G476));
  not1  g1037(.din(new_new_n981__), .dout(G477));
  not1  g1038(.din(new_new_n986__), .dout(G478));
  not1  g1039(.din(new_new_n991__), .dout(G479));
  not1  g1040(.din(new_new_n1004__), .dout(G480));
  not1  g1041(.din(new_new_n1009__), .dout(G481));
  not1  g1042(.din(new_new_n1014__), .dout(G482));
  not1  g1043(.din(new_new_n1019__), .dout(G483));
  not1  g1044(.din(new_new_n1032__), .dout(G484));
  not1  g1045(.din(new_new_n1037__), .dout(G485));
  not1  g1046(.din(new_new_n1042__), .dout(G486));
  not1  g1047(.din(new_new_n1047__), .dout(G487));
  not1  g1048(.din(new_new_n1060__), .dout(G488));
  not1  g1049(.din(new_new_n1065__), .dout(G489));
  not1  g1050(.din(new_new_n1070__), .dout(G490));
  not1  g1051(.din(new_new_n1075__), .dout(G491));
  not1  g1052(.din(new_new_n1088__), .dout(G492));
  not1  g1053(.din(new_new_n1093__), .dout(G493));
  not1  g1054(.din(new_new_n1098__), .dout(G494));
  not1  g1055(.din(new_new_n1103__), .dout(G495));
  not1  g1056(.din(new_new_n1116__), .dout(G496));
  not1  g1057(.din(new_new_n1121__), .dout(G497));
  not1  g1058(.din(new_new_n1126__), .dout(G498));
  not1  g1059(.din(new_new_n1131__), .dout(G499));
  not1  g1060(.din(new_new_n631__), .dout(n3791));
  not1  g1061(.din(new_new_n633__), .dout(n3794));
  not1  g1062(.din(new_new_n635__), .dout(n3797));
  not1  g1063(.din(new_new_n637__), .dout(n3800));
  not1  g1064(.din(new_new_n639__), .dout(n3803));
  not1  g1065(.din(new_new_n641__), .dout(n3806));
  not1  g1066(.din(new_new_n643__), .dout(n3809));
  not1  g1067(.din(new_new_n645__), .dout(n3812));
  not1  g1068(.din(new_new_n647__), .dout(n3815));
  not1  g1069(.din(new_new_n649__), .dout(n3818));
  not1  g1070(.din(new_new_n651__), .dout(n3821));
  not1  g1071(.din(new_new_n653__), .dout(n3824));
  not1  g1072(.din(new_new_n655__), .dout(n3827));
  not1  g1073(.din(new_new_n657__), .dout(n3830));
  not1  g1074(.din(new_new_n659__), .dout(n3833));
  not1  g1075(.din(new_new_n661__), .dout(n3836));
  not1  g1076(.din(new_new_n663__), .dout(n3839));
  not1  g1077(.din(new_new_n665__), .dout(n3842));
  not1  g1078(.din(new_new_n667__), .dout(n3845));
  not1  g1079(.din(new_new_n669__), .dout(n3848));
  not1  g1080(.din(new_new_n671__), .dout(n3851));
  not1  g1081(.din(new_new_n673__), .dout(n3854));
  not1  g1082(.din(new_new_n675__), .dout(n3857));
  not1  g1083(.din(new_new_n677__), .dout(n3860));
  not1  g1084(.din(new_new_n679__), .dout(n3863));
  not1  g1085(.din(new_new_n681__), .dout(n3866));
  not1  g1086(.din(new_new_n683__), .dout(n3869));
  not1  g1087(.din(new_new_n685__), .dout(n3872));
  not1  g1088(.din(new_new_n687__), .dout(n3875));
  not1  g1089(.din(new_new_n689__), .dout(n3878));
  not1  g1090(.din(new_new_n691__), .dout(n3881));
  not1  g1091(.din(new_new_n693__), .dout(n3884));
  not1  g1092(.din(new_new_n515__), .dout(n3887));
  not1  g1093(.din(new_new_n517__), .dout(n3890));
  not1  g1094(.din(new_new_n519__), .dout(n3893));
  not1  g1095(.din(new_new_n521__), .dout(n3896));
  not1  g1096(.din(new_new_n523__), .dout(n3899));
  not1  g1097(.din(new_new_n525__), .dout(n3902));
  not1  g1098(.din(new_new_n527__), .dout(n3905));
  not1  g1099(.din(new_new_n529__), .dout(n3908));
  not1  g1100(.din(new_new_n531__), .dout(n3911));
  not1  g1101(.din(new_new_n1937__), .dout(n3914));
  not1  g1102(.din(new_new_n1934__), .dout(n3917));
  not1  g1103(.din(new_new_n1929__), .dout(n3920));
  not1  g1104(.din(new_new_n1926__), .dout(n3923));
  not1  g1105(.din(new_new_n1956__), .dout(n3926));
  not1  g1106(.din(new_new_n1953__), .dout(n3929));
  not1  g1107(.din(new_new_n1948__), .dout(n3932));
  not1  g1108(.din(new_new_n1945__), .dout(n3935));
  not1  g1109(.din(new_new_n1959__), .dout(n3938));
  not1  g1110(.din(new_new_n2005__), .dout(n3941));
  not1  g1111(.din(new_new_n2037__), .dout(n3944));
  not1  g1112(.din(new_new_n2057__), .dout(n3947));
  not1  g1113(.din(new_new_n1961__), .dout(n3950));
  not1  g1114(.din(new_new_n2007__), .dout(n3953));
  not1  g1115(.din(new_new_n2039__), .dout(n3956));
  not1  g1116(.din(new_new_n2059__), .dout(n3959));
  not1  g1117(.din(new_new_n1965__), .dout(n3962));
  not1  g1118(.din(new_new_n2011__), .dout(n3965));
  not1  g1119(.din(new_new_n2043__), .dout(n3968));
  not1  g1120(.din(new_new_n2063__), .dout(n3971));
  not1  g1121(.din(new_new_n1967__), .dout(n3974));
  not1  g1122(.din(new_new_n2013__), .dout(n3977));
  not1  g1123(.din(new_new_n2045__), .dout(n3980));
  not1  g1124(.din(new_new_n2065__), .dout(n3983));
  not1  g1125(.din(new_new_n2077__), .dout(n3986));
  not1  g1126(.din(new_new_n2109__), .dout(n3989));
  not1  g1127(.din(new_new_n2141__), .dout(n3992));
  not1  g1128(.din(new_new_n2161__), .dout(n3995));
  not1  g1129(.din(new_new_n2079__), .dout(n3998));
  not1  g1130(.din(new_new_n2111__), .dout(n4001));
  not1  g1131(.din(new_new_n2143__), .dout(n4004));
  not1  g1132(.din(new_new_n2163__), .dout(n4007));
  not1  g1133(.din(new_new_n2083__), .dout(n4010));
  not1  g1134(.din(new_new_n2115__), .dout(n4013));
  not1  g1135(.din(new_new_n2147__), .dout(n4016));
  not1  g1136(.din(new_new_n2167__), .dout(n4019));
  not1  g1137(.din(new_new_n2085__), .dout(n4022));
  not1  g1138(.din(new_new_n2117__), .dout(n4025));
  not1  g1139(.din(new_new_n2149__), .dout(n4028));
  not1  g1140(.din(new_new_n2169__), .dout(n4031));
  not1  g1141(.din(new_new_n1938__), .dout(n4034));
  buf1  g1142(.din(n4034), .dout(n4037));
  not1  g1143(.din(new_new_n1935__), .dout(n4040));
  buf1  g1144(.din(n4040), .dout(n4043));
  not1  g1145(.din(new_new_n1930__), .dout(n4046));
  buf1  g1146(.din(n4046), .dout(n4049));
  not1  g1147(.din(new_new_n1927__), .dout(n4052));
  buf1  g1148(.din(n4052), .dout(n4055));
  not1  g1149(.din(new_new_n1957__), .dout(n4058));
  buf1  g1150(.din(n4058), .dout(n4061));
  not1  g1151(.din(new_new_n1954__), .dout(n4064));
  buf1  g1152(.din(n4064), .dout(n4067));
  not1  g1153(.din(new_new_n1949__), .dout(n4070));
  buf1  g1154(.din(n4070), .dout(n4073));
  not1  g1155(.din(new_new_n1946__), .dout(n4076));
  buf1  g1156(.din(n4076), .dout(n4079));
  not1  g1157(.din(new_new_n1145__), .dout(n4082));
  not1  g1158(.din(new_new_n1159__), .dout(n4085));
  not1  g1159(.din(new_new_n2181__), .dout(n4088));
  not1  g1160(.din(new_new_n2183__), .dout(n4091));
  not1  g1161(.din(new_new_n2187__), .dout(n4094));
  not1  g1162(.din(new_new_n2189__), .dout(n4097));
  not1  g1163(.din(new_new_n2193__), .dout(n4100));
  not1  g1164(.din(new_new_n2195__), .dout(n4103));
  not1  g1165(.din(new_new_n2199__), .dout(n4106));
  not1  g1166(.din(new_new_n2201__), .dout(n4109));
  not1  g1167(.din(new_new_n2205__), .dout(n4112));
  not1  g1168(.din(new_new_n2207__), .dout(n4115));
  not1  g1169(.din(new_new_n2211__), .dout(n4118));
  not1  g1170(.din(new_new_n2213__), .dout(n4121));
  not1  g1171(.din(new_new_n2217__), .dout(n4124));
  not1  g1172(.din(new_new_n2219__), .dout(n4127));
  not1  g1173(.din(new_new_n2223__), .dout(n4130));
  not1  g1174(.din(new_new_n2225__), .dout(n4133));
  not1  g1175(.din(new_new_n2229__), .dout(n4136));
  not1  g1176(.din(new_new_n2231__), .dout(n4139));
  not1  g1177(.din(new_new_n2235__), .dout(n4142));
  not1  g1178(.din(new_new_n2237__), .dout(n4145));
  not1  g1179(.din(new_new_n2241__), .dout(n4148));
  not1  g1180(.din(new_new_n2243__), .dout(n4151));
  not1  g1181(.din(new_new_n2247__), .dout(n4154));
  not1  g1182(.din(new_new_n2249__), .dout(n4157));
  not1  g1183(.din(new_new_n2253__), .dout(n4160));
  not1  g1184(.din(new_new_n2255__), .dout(n4163));
  not1  g1185(.din(new_new_n2259__), .dout(n4166));
  not1  g1186(.din(new_new_n2261__), .dout(n4169));
  not1  g1187(.din(new_new_n2265__), .dout(n4172));
  not1  g1188(.din(new_new_n2267__), .dout(n4175));
  not1  g1189(.din(new_new_n2271__), .dout(n4178));
  not1  g1190(.din(new_new_n2273__), .dout(n4181));
  not1  g1191(.din(new_new_n1194__), .dout(n4184));
  not1  g1192(.din(new_new_n1229__), .dout(n4187));
  not1  g1193(.din(new_new_n1264__), .dout(n4190));
  not1  g1194(.din(new_new_n1299__), .dout(n4193));
  not1  g1195(.din(new_new_n1334__), .dout(n4196));
  not1  g1196(.din(new_new_n1369__), .dout(n4199));
  not1  g1197(.din(new_new_n1404__), .dout(n4202));
  not1  g1198(.din(new_new_n1439__), .dout(n4205));
  not1  g1199(.din(new_new_n597__), .dout(n4208));
  not1  g1200(.din(new_new_n599__), .dout(n4211));
  not1  g1201(.din(new_new_n601__), .dout(n4214));
  not1  g1202(.din(new_new_n603__), .dout(n4217));
  not1  g1203(.din(new_new_n605__), .dout(n4220));
  not1  g1204(.din(new_new_n607__), .dout(n4223));
  not1  g1205(.din(new_new_n609__), .dout(n4226));
  not1  g1206(.din(new_new_n611__), .dout(n4229));
  not1  g1207(.din(new_new_n613__), .dout(n4232));
  not1  g1208(.din(new_new_n1454__), .dout(n4235));
  not1  g1209(.din(new_new_n1469__), .dout(n4238));
  not1  g1210(.din(new_new_n1484__), .dout(n4241));
  not1  g1211(.din(new_new_n1499__), .dout(n4244));
  not1  g1212(.din(new_new_n1514__), .dout(n4247));
  not1  g1213(.din(new_new_n1529__), .dout(n4250));
  not1  g1214(.din(new_new_n1544__), .dout(n4253));
  not1  g1215(.din(new_new_n1559__), .dout(n4256));
  not1  g1216(.din(new_new_n451__), .dout(n4259));
  not1  g1217(.din(new_new_n453__), .dout(n4262));
  not1  g1218(.din(new_new_n455__), .dout(n4265));
  not1  g1219(.din(new_new_n457__), .dout(n4268));
  not1  g1220(.din(new_new_n459__), .dout(n4271));
  not1  g1221(.din(new_new_n461__), .dout(n4274));
  not1  g1222(.din(new_new_n463__), .dout(n4277));
  not1  g1223(.din(new_new_n465__), .dout(n4280));
  not1  g1224(.din(new_new_n467__), .dout(n4283));
  not1  g1225(.din(new_new_n469__), .dout(n4286));
  not1  g1226(.din(new_new_n471__), .dout(n4289));
  not1  g1227(.din(new_new_n473__), .dout(n4292));
  not1  g1228(.din(new_new_n475__), .dout(n4295));
  not1  g1229(.din(new_new_n477__), .dout(n4298));
  not1  g1230(.din(new_new_n479__), .dout(n4301));
  not1  g1231(.din(new_new_n481__), .dout(n4304));
  not1  g1232(.din(new_new_n483__), .dout(n4307));
  not1  g1233(.din(new_new_n485__), .dout(n4310));
  not1  g1234(.din(new_new_n487__), .dout(n4313));
  not1  g1235(.din(new_new_n489__), .dout(n4316));
  not1  g1236(.din(new_new_n491__), .dout(n4319));
  not1  g1237(.din(new_new_n493__), .dout(n4322));
  not1  g1238(.din(new_new_n495__), .dout(n4325));
  not1  g1239(.din(new_new_n497__), .dout(n4328));
  not1  g1240(.din(new_new_n499__), .dout(n4331));
  not1  g1241(.din(new_new_n501__), .dout(n4334));
  not1  g1242(.din(new_new_n503__), .dout(n4337));
  not1  g1243(.din(new_new_n505__), .dout(n4340));
  not1  g1244(.din(new_new_n507__), .dout(n4343));
  not1  g1245(.din(new_new_n509__), .dout(n4346));
  not1  g1246(.din(new_new_n511__), .dout(n4349));
  not1  g1247(.din(new_new_n513__), .dout(n4352));
  buf1  g1248(.din(new_new_n622__), .dout(new_new_n1780__));
  buf1  g1249(.din(new_new_n1780__), .dout(new_new_n1781__));
  buf1  g1250(.din(new_new_n1781__), .dout(new_new_n1782__));
  buf1  g1251(.din(new_new_n1781__), .dout(new_new_n1783__));
  buf1  g1252(.din(new_new_n1780__), .dout(new_new_n1784__));
  buf1  g1253(.din(new_new_n623__), .dout(new_new_n1785__));
  buf1  g1254(.din(new_new_n1785__), .dout(new_new_n1786__));
  buf1  g1255(.din(new_new_n1786__), .dout(new_new_n1787__));
  buf1  g1256(.din(new_new_n1786__), .dout(new_new_n1788__));
  buf1  g1257(.din(new_new_n1785__), .dout(new_new_n1789__));
  buf1  g1258(.din(new_new_n626__), .dout(new_new_n1790__));
  buf1  g1259(.din(new_new_n1790__), .dout(new_new_n1791__));
  buf1  g1260(.din(new_new_n1791__), .dout(new_new_n1792__));
  buf1  g1261(.din(new_new_n1791__), .dout(new_new_n1793__));
  buf1  g1262(.din(new_new_n1790__), .dout(new_new_n1794__));
  buf1  g1263(.din(new_new_n627__), .dout(new_new_n1795__));
  buf1  g1264(.din(new_new_n1795__), .dout(new_new_n1796__));
  buf1  g1265(.din(new_new_n1796__), .dout(new_new_n1797__));
  buf1  g1266(.din(new_new_n1796__), .dout(new_new_n1798__));
  buf1  g1267(.din(new_new_n1795__), .dout(new_new_n1799__));
  buf1  g1268(.din(new_new_n726__), .dout(new_new_n1800__));
  buf1  g1269(.din(new_new_n1800__), .dout(new_new_n1801__));
  buf1  g1270(.din(new_new_n1800__), .dout(new_new_n1802__));
  buf1  g1271(.din(new_new_n727__), .dout(new_new_n1803__));
  buf1  g1272(.din(new_new_n1803__), .dout(new_new_n1804__));
  buf1  g1273(.din(new_new_n1803__), .dout(new_new_n1805__));
  buf1  g1274(.din(new_new_n914__), .dout(new_new_n1806__));
  buf1  g1275(.din(new_new_n1806__), .dout(new_new_n1807__));
  buf1  g1276(.din(new_new_n1806__), .dout(new_new_n1808__));
  buf1  g1277(.din(new_new_n614__), .dout(new_new_n1809__));
  buf1  g1278(.din(new_new_n1809__), .dout(new_new_n1810__));
  buf1  g1279(.din(new_new_n1810__), .dout(new_new_n1811__));
  buf1  g1280(.din(new_new_n1810__), .dout(new_new_n1812__));
  buf1  g1281(.din(new_new_n1809__), .dout(new_new_n1813__));
  buf1  g1282(.din(new_new_n915__), .dout(new_new_n1814__));
  buf1  g1283(.din(new_new_n1814__), .dout(new_new_n1815__));
  buf1  g1284(.din(new_new_n1814__), .dout(new_new_n1816__));
  buf1  g1285(.din(new_new_n615__), .dout(new_new_n1817__));
  buf1  g1286(.din(new_new_n1817__), .dout(new_new_n1818__));
  buf1  g1287(.din(new_new_n1818__), .dout(new_new_n1819__));
  buf1  g1288(.din(new_new_n1818__), .dout(new_new_n1820__));
  buf1  g1289(.din(new_new_n1817__), .dout(new_new_n1821__));
  buf1  g1290(.din(new_new_n616__), .dout(new_new_n1822__));
  buf1  g1291(.din(new_new_n1822__), .dout(new_new_n1823__));
  buf1  g1292(.din(new_new_n1823__), .dout(new_new_n1824__));
  buf1  g1293(.din(new_new_n1823__), .dout(new_new_n1825__));
  buf1  g1294(.din(new_new_n1822__), .dout(new_new_n1826__));
  buf1  g1295(.din(new_new_n617__), .dout(new_new_n1827__));
  buf1  g1296(.din(new_new_n1827__), .dout(new_new_n1828__));
  buf1  g1297(.din(new_new_n1828__), .dout(new_new_n1829__));
  buf1  g1298(.din(new_new_n1828__), .dout(new_new_n1830__));
  buf1  g1299(.din(new_new_n1827__), .dout(new_new_n1831__));
  buf1  g1300(.din(new_new_n618__), .dout(new_new_n1832__));
  buf1  g1301(.din(new_new_n1832__), .dout(new_new_n1833__));
  buf1  g1302(.din(new_new_n1833__), .dout(new_new_n1834__));
  buf1  g1303(.din(new_new_n1833__), .dout(new_new_n1835__));
  buf1  g1304(.din(new_new_n1832__), .dout(new_new_n1836__));
  buf1  g1305(.din(new_new_n619__), .dout(new_new_n1837__));
  buf1  g1306(.din(new_new_n1837__), .dout(new_new_n1838__));
  buf1  g1307(.din(new_new_n1838__), .dout(new_new_n1839__));
  buf1  g1308(.din(new_new_n1838__), .dout(new_new_n1840__));
  buf1  g1309(.din(new_new_n1837__), .dout(new_new_n1841__));
  buf1  g1310(.din(new_new_n620__), .dout(new_new_n1842__));
  buf1  g1311(.din(new_new_n1842__), .dout(new_new_n1843__));
  buf1  g1312(.din(new_new_n1843__), .dout(new_new_n1844__));
  buf1  g1313(.din(new_new_n1843__), .dout(new_new_n1845__));
  buf1  g1314(.din(new_new_n1842__), .dout(new_new_n1846__));
  buf1  g1315(.din(new_new_n621__), .dout(new_new_n1847__));
  buf1  g1316(.din(new_new_n1847__), .dout(new_new_n1848__));
  buf1  g1317(.din(new_new_n1848__), .dout(new_new_n1849__));
  buf1  g1318(.din(new_new_n1848__), .dout(new_new_n1850__));
  buf1  g1319(.din(new_new_n1847__), .dout(new_new_n1851__));
  buf1  g1320(.din(new_new_n628__), .dout(new_new_n1852__));
  buf1  g1321(.din(new_new_n1852__), .dout(new_new_n1853__));
  buf1  g1322(.din(new_new_n1853__), .dout(new_new_n1854__));
  buf1  g1323(.din(new_new_n1853__), .dout(new_new_n1855__));
  buf1  g1324(.din(new_new_n1852__), .dout(new_new_n1856__));
  buf1  g1325(.din(new_new_n629__), .dout(new_new_n1857__));
  buf1  g1326(.din(new_new_n1857__), .dout(new_new_n1858__));
  buf1  g1327(.din(new_new_n1858__), .dout(new_new_n1859__));
  buf1  g1328(.din(new_new_n1858__), .dout(new_new_n1860__));
  buf1  g1329(.din(new_new_n1857__), .dout(new_new_n1861__));
  buf1  g1330(.din(new_new_n942__), .dout(new_new_n1862__));
  buf1  g1331(.din(new_new_n1862__), .dout(new_new_n1863__));
  buf1  g1332(.din(new_new_n1862__), .dout(new_new_n1864__));
  buf1  g1333(.din(new_new_n943__), .dout(new_new_n1865__));
  buf1  g1334(.din(new_new_n1865__), .dout(new_new_n1866__));
  buf1  g1335(.din(new_new_n1865__), .dout(new_new_n1867__));
  buf1  g1336(.din(new_new_n624__), .dout(new_new_n1868__));
  buf1  g1337(.din(new_new_n1868__), .dout(new_new_n1869__));
  buf1  g1338(.din(new_new_n1869__), .dout(new_new_n1870__));
  buf1  g1339(.din(new_new_n1869__), .dout(new_new_n1871__));
  buf1  g1340(.din(new_new_n1868__), .dout(new_new_n1872__));
  buf1  g1341(.din(new_new_n625__), .dout(new_new_n1873__));
  buf1  g1342(.din(new_new_n1873__), .dout(new_new_n1874__));
  buf1  g1343(.din(new_new_n1874__), .dout(new_new_n1875__));
  buf1  g1344(.din(new_new_n1874__), .dout(new_new_n1876__));
  buf1  g1345(.din(new_new_n1873__), .dout(new_new_n1877__));
  buf1  g1346(.din(new_new_n970__), .dout(new_new_n1878__));
  buf1  g1347(.din(new_new_n1878__), .dout(new_new_n1879__));
  buf1  g1348(.din(new_new_n1878__), .dout(new_new_n1880__));
  buf1  g1349(.din(new_new_n971__), .dout(new_new_n1881__));
  buf1  g1350(.din(new_new_n1881__), .dout(new_new_n1882__));
  buf1  g1351(.din(new_new_n1881__), .dout(new_new_n1883__));
  buf1  g1352(.din(new_new_n998__), .dout(new_new_n1884__));
  buf1  g1353(.din(new_new_n1884__), .dout(new_new_n1885__));
  buf1  g1354(.din(new_new_n1884__), .dout(new_new_n1886__));
  buf1  g1355(.din(new_new_n999__), .dout(new_new_n1887__));
  buf1  g1356(.din(new_new_n1887__), .dout(new_new_n1888__));
  buf1  g1357(.din(new_new_n1887__), .dout(new_new_n1889__));
  buf1  g1358(.din(new_new_n728__), .dout(new_new_n1890__));
  buf1  g1359(.din(new_new_n1890__), .dout(new_new_n1891__));
  buf1  g1360(.din(new_new_n1890__), .dout(new_new_n1892__));
  buf1  g1361(.din(new_new_n729__), .dout(new_new_n1893__));
  buf1  g1362(.din(new_new_n1893__), .dout(new_new_n1894__));
  buf1  g1363(.din(new_new_n1893__), .dout(new_new_n1895__));
  buf1  g1364(.din(new_new_n1026__), .dout(new_new_n1896__));
  buf1  g1365(.din(new_new_n1896__), .dout(new_new_n1897__));
  buf1  g1366(.din(new_new_n1896__), .dout(new_new_n1898__));
  buf1  g1367(.din(new_new_n1027__), .dout(new_new_n1899__));
  buf1  g1368(.din(new_new_n1899__), .dout(new_new_n1900__));
  buf1  g1369(.din(new_new_n1899__), .dout(new_new_n1901__));
  buf1  g1370(.din(new_new_n1054__), .dout(new_new_n1902__));
  buf1  g1371(.din(new_new_n1902__), .dout(new_new_n1903__));
  buf1  g1372(.din(new_new_n1902__), .dout(new_new_n1904__));
  buf1  g1373(.din(new_new_n1055__), .dout(new_new_n1905__));
  buf1  g1374(.din(new_new_n1905__), .dout(new_new_n1906__));
  buf1  g1375(.din(new_new_n1905__), .dout(new_new_n1907__));
  buf1  g1376(.din(new_new_n1082__), .dout(new_new_n1908__));
  buf1  g1377(.din(new_new_n1908__), .dout(new_new_n1909__));
  buf1  g1378(.din(new_new_n1908__), .dout(new_new_n1910__));
  buf1  g1379(.din(new_new_n1083__), .dout(new_new_n1911__));
  buf1  g1380(.din(new_new_n1911__), .dout(new_new_n1912__));
  buf1  g1381(.din(new_new_n1911__), .dout(new_new_n1913__));
  buf1  g1382(.din(new_new_n1110__), .dout(new_new_n1914__));
  buf1  g1383(.din(new_new_n1914__), .dout(new_new_n1915__));
  buf1  g1384(.din(new_new_n1914__), .dout(new_new_n1916__));
  buf1  g1385(.din(new_new_n1111__), .dout(new_new_n1917__));
  buf1  g1386(.din(new_new_n1917__), .dout(new_new_n1918__));
  buf1  g1387(.din(new_new_n1917__), .dout(new_new_n1919__));
  buf1  g1388(.din(new_new_n796__), .dout(new_new_n1920__));
  buf1  g1389(.din(new_new_n794__), .dout(new_new_n1921__));
  buf1  g1390(.din(new_new_n1132__), .dout(new_new_n1922__));
  buf1  g1391(.din(new_new_n798__), .dout(new_new_n1923__));
  buf1  g1392(.din(new_new_n1923__), .dout(new_new_n1924__));
  buf1  g1393(.din(new_new_n801__), .dout(new_new_n1925__));
  buf1  g1394(.din(new_new_n1925__), .dout(new_new_n1926__));
  buf1  g1395(.din(new_new_n1925__), .dout(new_new_n1927__));
  buf1  g1396(.din(new_new_n799__), .dout(new_new_n1928__));
  buf1  g1397(.din(new_new_n1928__), .dout(new_new_n1929__));
  buf1  g1398(.din(new_new_n1928__), .dout(new_new_n1930__));
  buf1  g1399(.din(new_new_n800__), .dout(new_new_n1931__));
  buf1  g1400(.din(new_new_n1931__), .dout(new_new_n1932__));
  buf1  g1401(.din(new_new_n797__), .dout(new_new_n1933__));
  buf1  g1402(.din(new_new_n1933__), .dout(new_new_n1934__));
  buf1  g1403(.din(new_new_n1933__), .dout(new_new_n1935__));
  buf1  g1404(.din(new_new_n795__), .dout(new_new_n1936__));
  buf1  g1405(.din(new_new_n1936__), .dout(new_new_n1937__));
  buf1  g1406(.din(new_new_n1936__), .dout(new_new_n1938__));
  buf1  g1407(.din(new_new_n804__), .dout(new_new_n1939__));
  buf1  g1408(.din(new_new_n802__), .dout(new_new_n1940__));
  buf1  g1409(.din(new_new_n1146__), .dout(new_new_n1941__));
  buf1  g1410(.din(new_new_n806__), .dout(new_new_n1942__));
  buf1  g1411(.din(new_new_n1942__), .dout(new_new_n1943__));
  buf1  g1412(.din(new_new_n809__), .dout(new_new_n1944__));
  buf1  g1413(.din(new_new_n1944__), .dout(new_new_n1945__));
  buf1  g1414(.din(new_new_n1944__), .dout(new_new_n1946__));
  buf1  g1415(.din(new_new_n807__), .dout(new_new_n1947__));
  buf1  g1416(.din(new_new_n1947__), .dout(new_new_n1948__));
  buf1  g1417(.din(new_new_n1947__), .dout(new_new_n1949__));
  buf1  g1418(.din(new_new_n808__), .dout(new_new_n1950__));
  buf1  g1419(.din(new_new_n1950__), .dout(new_new_n1951__));
  buf1  g1420(.din(new_new_n805__), .dout(new_new_n1952__));
  buf1  g1421(.din(new_new_n1952__), .dout(new_new_n1953__));
  buf1  g1422(.din(new_new_n1952__), .dout(new_new_n1954__));
  buf1  g1423(.din(new_new_n803__), .dout(new_new_n1955__));
  buf1  g1424(.din(new_new_n1955__), .dout(new_new_n1956__));
  buf1  g1425(.din(new_new_n1955__), .dout(new_new_n1957__));
  buf1  g1426(.din(new_new_n738__), .dout(new_new_n1958__));
  buf1  g1427(.din(new_new_n731__), .dout(new_new_n1959__));
  buf1  g1428(.din(new_new_n1959__), .dout(new_new_n1960__));
  buf1  g1429(.din(new_new_n739__), .dout(new_new_n1961__));
  buf1  g1430(.din(new_new_n1961__), .dout(new_new_n1962__));
  buf1  g1431(.din(new_new_n730__), .dout(new_new_n1963__));
  buf1  g1432(.din(new_new_n754__), .dout(new_new_n1964__));
  buf1  g1433(.din(new_new_n747__), .dout(new_new_n1965__));
  buf1  g1434(.din(new_new_n1965__), .dout(new_new_n1966__));
  buf1  g1435(.din(new_new_n755__), .dout(new_new_n1967__));
  buf1  g1436(.din(new_new_n1967__), .dout(new_new_n1968__));
  buf1  g1437(.din(new_new_n746__), .dout(new_new_n1969__));
  buf1  g1438(.din(new_new_n1171__), .dout(new_new_n1970__));
  buf1  g1439(.din(new_new_n1164__), .dout(new_new_n1971__));
  buf1  g1440(.din(new_new_n1170__), .dout(new_new_n1972__));
  buf1  g1441(.din(new_new_n1165__), .dout(new_new_n1973__));
  buf1  g1442(.din(new_new_n826__), .dout(new_new_n1974__));
  buf1  g1443(.din(new_new_n1974__), .dout(new_new_n1975__));
  buf1  g1444(.din(new_new_n1975__), .dout(new_new_n1976__));
  buf1  g1445(.din(new_new_n1975__), .dout(new_new_n1977__));
  buf1  g1446(.din(new_new_n1974__), .dout(new_new_n1978__));
  buf1  g1447(.din(new_new_n1978__), .dout(new_new_n1979__));
  buf1  g1448(.din(new_new_n1978__), .dout(new_new_n1980__));
  buf1  g1449(.din(new_new_n827__), .dout(new_new_n1981__));
  buf1  g1450(.din(new_new_n1981__), .dout(new_new_n1982__));
  buf1  g1451(.din(new_new_n1982__), .dout(new_new_n1983__));
  buf1  g1452(.din(new_new_n1982__), .dout(new_new_n1984__));
  buf1  g1453(.din(new_new_n1981__), .dout(new_new_n1985__));
  buf1  g1454(.din(new_new_n1985__), .dout(new_new_n1986__));
  buf1  g1455(.din(new_new_n1985__), .dout(new_new_n1987__));
  buf1  g1456(.din(new_new_n838__), .dout(new_new_n1988__));
  buf1  g1457(.din(new_new_n1988__), .dout(new_new_n1989__));
  buf1  g1458(.din(new_new_n1988__), .dout(new_new_n1990__));
  buf1  g1459(.din(new_new_n837__), .dout(new_new_n1991__));
  buf1  g1460(.din(new_new_n1991__), .dout(new_new_n1992__));
  buf1  g1461(.din(new_new_n1991__), .dout(new_new_n1993__));
  buf1  g1462(.din(new_new_n839__), .dout(new_new_n1994__));
  buf1  g1463(.din(new_new_n1994__), .dout(new_new_n1995__));
  buf1  g1464(.din(new_new_n1994__), .dout(new_new_n1996__));
  buf1  g1465(.din(new_new_n836__), .dout(new_new_n1997__));
  buf1  g1466(.din(new_new_n1997__), .dout(new_new_n1998__));
  buf1  g1467(.din(new_new_n1997__), .dout(new_new_n1999__));
  buf1  g1468(.din(new_new_n1185__), .dout(new_new_n2000__));
  buf1  g1469(.din(new_new_n1179__), .dout(new_new_n2001__));
  buf1  g1470(.din(new_new_n1184__), .dout(new_new_n2002__));
  buf1  g1471(.din(new_new_n1178__), .dout(new_new_n2003__));
  buf1  g1472(.din(new_new_n740__), .dout(new_new_n2004__));
  buf1  g1473(.din(new_new_n733__), .dout(new_new_n2005__));
  buf1  g1474(.din(new_new_n2005__), .dout(new_new_n2006__));
  buf1  g1475(.din(new_new_n741__), .dout(new_new_n2007__));
  buf1  g1476(.din(new_new_n2007__), .dout(new_new_n2008__));
  buf1  g1477(.din(new_new_n732__), .dout(new_new_n2009__));
  buf1  g1478(.din(new_new_n756__), .dout(new_new_n2010__));
  buf1  g1479(.din(new_new_n749__), .dout(new_new_n2011__));
  buf1  g1480(.din(new_new_n2011__), .dout(new_new_n2012__));
  buf1  g1481(.din(new_new_n757__), .dout(new_new_n2013__));
  buf1  g1482(.din(new_new_n2013__), .dout(new_new_n2014__));
  buf1  g1483(.din(new_new_n748__), .dout(new_new_n2015__));
  buf1  g1484(.din(new_new_n1206__), .dout(new_new_n2016__));
  buf1  g1485(.din(new_new_n1199__), .dout(new_new_n2017__));
  buf1  g1486(.din(new_new_n1205__), .dout(new_new_n2018__));
  buf1  g1487(.din(new_new_n1200__), .dout(new_new_n2019__));
  buf1  g1488(.din(new_new_n842__), .dout(new_new_n2020__));
  buf1  g1489(.din(new_new_n2020__), .dout(new_new_n2021__));
  buf1  g1490(.din(new_new_n2020__), .dout(new_new_n2022__));
  buf1  g1491(.din(new_new_n841__), .dout(new_new_n2023__));
  buf1  g1492(.din(new_new_n2023__), .dout(new_new_n2024__));
  buf1  g1493(.din(new_new_n2023__), .dout(new_new_n2025__));
  buf1  g1494(.din(new_new_n843__), .dout(new_new_n2026__));
  buf1  g1495(.din(new_new_n2026__), .dout(new_new_n2027__));
  buf1  g1496(.din(new_new_n2026__), .dout(new_new_n2028__));
  buf1  g1497(.din(new_new_n840__), .dout(new_new_n2029__));
  buf1  g1498(.din(new_new_n2029__), .dout(new_new_n2030__));
  buf1  g1499(.din(new_new_n2029__), .dout(new_new_n2031__));
  buf1  g1500(.din(new_new_n1220__), .dout(new_new_n2032__));
  buf1  g1501(.din(new_new_n1214__), .dout(new_new_n2033__));
  buf1  g1502(.din(new_new_n1219__), .dout(new_new_n2034__));
  buf1  g1503(.din(new_new_n1213__), .dout(new_new_n2035__));
  buf1  g1504(.din(new_new_n742__), .dout(new_new_n2036__));
  buf1  g1505(.din(new_new_n735__), .dout(new_new_n2037__));
  buf1  g1506(.din(new_new_n2037__), .dout(new_new_n2038__));
  buf1  g1507(.din(new_new_n743__), .dout(new_new_n2039__));
  buf1  g1508(.din(new_new_n2039__), .dout(new_new_n2040__));
  buf1  g1509(.din(new_new_n734__), .dout(new_new_n2041__));
  buf1  g1510(.din(new_new_n758__), .dout(new_new_n2042__));
  buf1  g1511(.din(new_new_n751__), .dout(new_new_n2043__));
  buf1  g1512(.din(new_new_n2043__), .dout(new_new_n2044__));
  buf1  g1513(.din(new_new_n759__), .dout(new_new_n2045__));
  buf1  g1514(.din(new_new_n2045__), .dout(new_new_n2046__));
  buf1  g1515(.din(new_new_n750__), .dout(new_new_n2047__));
  buf1  g1516(.din(new_new_n1241__), .dout(new_new_n2048__));
  buf1  g1517(.din(new_new_n1234__), .dout(new_new_n2049__));
  buf1  g1518(.din(new_new_n1240__), .dout(new_new_n2050__));
  buf1  g1519(.din(new_new_n1235__), .dout(new_new_n2051__));
  buf1  g1520(.din(new_new_n1255__), .dout(new_new_n2052__));
  buf1  g1521(.din(new_new_n1249__), .dout(new_new_n2053__));
  buf1  g1522(.din(new_new_n1254__), .dout(new_new_n2054__));
  buf1  g1523(.din(new_new_n1248__), .dout(new_new_n2055__));
  buf1  g1524(.din(new_new_n744__), .dout(new_new_n2056__));
  buf1  g1525(.din(new_new_n737__), .dout(new_new_n2057__));
  buf1  g1526(.din(new_new_n2057__), .dout(new_new_n2058__));
  buf1  g1527(.din(new_new_n745__), .dout(new_new_n2059__));
  buf1  g1528(.din(new_new_n2059__), .dout(new_new_n2060__));
  buf1  g1529(.din(new_new_n736__), .dout(new_new_n2061__));
  buf1  g1530(.din(new_new_n760__), .dout(new_new_n2062__));
  buf1  g1531(.din(new_new_n753__), .dout(new_new_n2063__));
  buf1  g1532(.din(new_new_n2063__), .dout(new_new_n2064__));
  buf1  g1533(.din(new_new_n761__), .dout(new_new_n2065__));
  buf1  g1534(.din(new_new_n2065__), .dout(new_new_n2066__));
  buf1  g1535(.din(new_new_n752__), .dout(new_new_n2067__));
  buf1  g1536(.din(new_new_n1276__), .dout(new_new_n2068__));
  buf1  g1537(.din(new_new_n1269__), .dout(new_new_n2069__));
  buf1  g1538(.din(new_new_n1275__), .dout(new_new_n2070__));
  buf1  g1539(.din(new_new_n1270__), .dout(new_new_n2071__));
  buf1  g1540(.din(new_new_n1290__), .dout(new_new_n2072__));
  buf1  g1541(.din(new_new_n1284__), .dout(new_new_n2073__));
  buf1  g1542(.din(new_new_n1289__), .dout(new_new_n2074__));
  buf1  g1543(.din(new_new_n1283__), .dout(new_new_n2075__));
  buf1  g1544(.din(new_new_n770__), .dout(new_new_n2076__));
  buf1  g1545(.din(new_new_n763__), .dout(new_new_n2077__));
  buf1  g1546(.din(new_new_n2077__), .dout(new_new_n2078__));
  buf1  g1547(.din(new_new_n771__), .dout(new_new_n2079__));
  buf1  g1548(.din(new_new_n2079__), .dout(new_new_n2080__));
  buf1  g1549(.din(new_new_n762__), .dout(new_new_n2081__));
  buf1  g1550(.din(new_new_n786__), .dout(new_new_n2082__));
  buf1  g1551(.din(new_new_n779__), .dout(new_new_n2083__));
  buf1  g1552(.din(new_new_n2083__), .dout(new_new_n2084__));
  buf1  g1553(.din(new_new_n787__), .dout(new_new_n2085__));
  buf1  g1554(.din(new_new_n2085__), .dout(new_new_n2086__));
  buf1  g1555(.din(new_new_n778__), .dout(new_new_n2087__));
  buf1  g1556(.din(new_new_n1311__), .dout(new_new_n2088__));
  buf1  g1557(.din(new_new_n1304__), .dout(new_new_n2089__));
  buf1  g1558(.din(new_new_n1310__), .dout(new_new_n2090__));
  buf1  g1559(.din(new_new_n1305__), .dout(new_new_n2091__));
  buf1  g1560(.din(new_new_n830__), .dout(new_new_n2092__));
  buf1  g1561(.din(new_new_n2092__), .dout(new_new_n2093__));
  buf1  g1562(.din(new_new_n2092__), .dout(new_new_n2094__));
  buf1  g1563(.din(new_new_n829__), .dout(new_new_n2095__));
  buf1  g1564(.din(new_new_n2095__), .dout(new_new_n2096__));
  buf1  g1565(.din(new_new_n2095__), .dout(new_new_n2097__));
  buf1  g1566(.din(new_new_n831__), .dout(new_new_n2098__));
  buf1  g1567(.din(new_new_n2098__), .dout(new_new_n2099__));
  buf1  g1568(.din(new_new_n2098__), .dout(new_new_n2100__));
  buf1  g1569(.din(new_new_n828__), .dout(new_new_n2101__));
  buf1  g1570(.din(new_new_n2101__), .dout(new_new_n2102__));
  buf1  g1571(.din(new_new_n2101__), .dout(new_new_n2103__));
  buf1  g1572(.din(new_new_n1325__), .dout(new_new_n2104__));
  buf1  g1573(.din(new_new_n1319__), .dout(new_new_n2105__));
  buf1  g1574(.din(new_new_n1324__), .dout(new_new_n2106__));
  buf1  g1575(.din(new_new_n1318__), .dout(new_new_n2107__));
  buf1  g1576(.din(new_new_n772__), .dout(new_new_n2108__));
  buf1  g1577(.din(new_new_n765__), .dout(new_new_n2109__));
  buf1  g1578(.din(new_new_n2109__), .dout(new_new_n2110__));
  buf1  g1579(.din(new_new_n773__), .dout(new_new_n2111__));
  buf1  g1580(.din(new_new_n2111__), .dout(new_new_n2112__));
  buf1  g1581(.din(new_new_n764__), .dout(new_new_n2113__));
  buf1  g1582(.din(new_new_n788__), .dout(new_new_n2114__));
  buf1  g1583(.din(new_new_n781__), .dout(new_new_n2115__));
  buf1  g1584(.din(new_new_n2115__), .dout(new_new_n2116__));
  buf1  g1585(.din(new_new_n789__), .dout(new_new_n2117__));
  buf1  g1586(.din(new_new_n2117__), .dout(new_new_n2118__));
  buf1  g1587(.din(new_new_n780__), .dout(new_new_n2119__));
  buf1  g1588(.din(new_new_n1346__), .dout(new_new_n2120__));
  buf1  g1589(.din(new_new_n1339__), .dout(new_new_n2121__));
  buf1  g1590(.din(new_new_n1345__), .dout(new_new_n2122__));
  buf1  g1591(.din(new_new_n1340__), .dout(new_new_n2123__));
  buf1  g1592(.din(new_new_n834__), .dout(new_new_n2124__));
  buf1  g1593(.din(new_new_n2124__), .dout(new_new_n2125__));
  buf1  g1594(.din(new_new_n2124__), .dout(new_new_n2126__));
  buf1  g1595(.din(new_new_n833__), .dout(new_new_n2127__));
  buf1  g1596(.din(new_new_n2127__), .dout(new_new_n2128__));
  buf1  g1597(.din(new_new_n2127__), .dout(new_new_n2129__));
  buf1  g1598(.din(new_new_n835__), .dout(new_new_n2130__));
  buf1  g1599(.din(new_new_n2130__), .dout(new_new_n2131__));
  buf1  g1600(.din(new_new_n2130__), .dout(new_new_n2132__));
  buf1  g1601(.din(new_new_n832__), .dout(new_new_n2133__));
  buf1  g1602(.din(new_new_n2133__), .dout(new_new_n2134__));
  buf1  g1603(.din(new_new_n2133__), .dout(new_new_n2135__));
  buf1  g1604(.din(new_new_n1360__), .dout(new_new_n2136__));
  buf1  g1605(.din(new_new_n1354__), .dout(new_new_n2137__));
  buf1  g1606(.din(new_new_n1359__), .dout(new_new_n2138__));
  buf1  g1607(.din(new_new_n1353__), .dout(new_new_n2139__));
  buf1  g1608(.din(new_new_n774__), .dout(new_new_n2140__));
  buf1  g1609(.din(new_new_n767__), .dout(new_new_n2141__));
  buf1  g1610(.din(new_new_n2141__), .dout(new_new_n2142__));
  buf1  g1611(.din(new_new_n775__), .dout(new_new_n2143__));
  buf1  g1612(.din(new_new_n2143__), .dout(new_new_n2144__));
  buf1  g1613(.din(new_new_n766__), .dout(new_new_n2145__));
  buf1  g1614(.din(new_new_n790__), .dout(new_new_n2146__));
  buf1  g1615(.din(new_new_n783__), .dout(new_new_n2147__));
  buf1  g1616(.din(new_new_n2147__), .dout(new_new_n2148__));
  buf1  g1617(.din(new_new_n791__), .dout(new_new_n2149__));
  buf1  g1618(.din(new_new_n2149__), .dout(new_new_n2150__));
  buf1  g1619(.din(new_new_n782__), .dout(new_new_n2151__));
  buf1  g1620(.din(new_new_n1381__), .dout(new_new_n2152__));
  buf1  g1621(.din(new_new_n1374__), .dout(new_new_n2153__));
  buf1  g1622(.din(new_new_n1380__), .dout(new_new_n2154__));
  buf1  g1623(.din(new_new_n1375__), .dout(new_new_n2155__));
  buf1  g1624(.din(new_new_n1395__), .dout(new_new_n2156__));
  buf1  g1625(.din(new_new_n1389__), .dout(new_new_n2157__));
  buf1  g1626(.din(new_new_n1394__), .dout(new_new_n2158__));
  buf1  g1627(.din(new_new_n1388__), .dout(new_new_n2159__));
  buf1  g1628(.din(new_new_n776__), .dout(new_new_n2160__));
  buf1  g1629(.din(new_new_n769__), .dout(new_new_n2161__));
  buf1  g1630(.din(new_new_n2161__), .dout(new_new_n2162__));
  buf1  g1631(.din(new_new_n777__), .dout(new_new_n2163__));
  buf1  g1632(.din(new_new_n2163__), .dout(new_new_n2164__));
  buf1  g1633(.din(new_new_n768__), .dout(new_new_n2165__));
  buf1  g1634(.din(new_new_n792__), .dout(new_new_n2166__));
  buf1  g1635(.din(new_new_n785__), .dout(new_new_n2167__));
  buf1  g1636(.din(new_new_n2167__), .dout(new_new_n2168__));
  buf1  g1637(.din(new_new_n793__), .dout(new_new_n2169__));
  buf1  g1638(.din(new_new_n2169__), .dout(new_new_n2170__));
  buf1  g1639(.din(new_new_n784__), .dout(new_new_n2171__));
  buf1  g1640(.din(new_new_n1416__), .dout(new_new_n2172__));
  buf1  g1641(.din(new_new_n1409__), .dout(new_new_n2173__));
  buf1  g1642(.din(new_new_n1415__), .dout(new_new_n2174__));
  buf1  g1643(.din(new_new_n1410__), .dout(new_new_n2175__));
  buf1  g1644(.din(new_new_n1430__), .dout(new_new_n2176__));
  buf1  g1645(.din(new_new_n1424__), .dout(new_new_n2177__));
  buf1  g1646(.din(new_new_n1429__), .dout(new_new_n2178__));
  buf1  g1647(.din(new_new_n1423__), .dout(new_new_n2179__));
  buf1  g1648(.din(new_new_n846__), .dout(new_new_n2180__));
  buf1  g1649(.din(new_new_n845__), .dout(new_new_n2181__));
  buf1  g1650(.din(new_new_n2181__), .dout(new_new_n2182__));
  buf1  g1651(.din(new_new_n847__), .dout(new_new_n2183__));
  buf1  g1652(.din(new_new_n2183__), .dout(new_new_n2184__));
  buf1  g1653(.din(new_new_n844__), .dout(new_new_n2185__));
  buf1  g1654(.din(new_new_n850__), .dout(new_new_n2186__));
  buf1  g1655(.din(new_new_n849__), .dout(new_new_n2187__));
  buf1  g1656(.din(new_new_n2187__), .dout(new_new_n2188__));
  buf1  g1657(.din(new_new_n851__), .dout(new_new_n2189__));
  buf1  g1658(.din(new_new_n2189__), .dout(new_new_n2190__));
  buf1  g1659(.din(new_new_n848__), .dout(new_new_n2191__));
  buf1  g1660(.din(new_new_n854__), .dout(new_new_n2192__));
  buf1  g1661(.din(new_new_n853__), .dout(new_new_n2193__));
  buf1  g1662(.din(new_new_n2193__), .dout(new_new_n2194__));
  buf1  g1663(.din(new_new_n855__), .dout(new_new_n2195__));
  buf1  g1664(.din(new_new_n2195__), .dout(new_new_n2196__));
  buf1  g1665(.din(new_new_n852__), .dout(new_new_n2197__));
  buf1  g1666(.din(new_new_n858__), .dout(new_new_n2198__));
  buf1  g1667(.din(new_new_n857__), .dout(new_new_n2199__));
  buf1  g1668(.din(new_new_n2199__), .dout(new_new_n2200__));
  buf1  g1669(.din(new_new_n859__), .dout(new_new_n2201__));
  buf1  g1670(.din(new_new_n2201__), .dout(new_new_n2202__));
  buf1  g1671(.din(new_new_n856__), .dout(new_new_n2203__));
  buf1  g1672(.din(new_new_n862__), .dout(new_new_n2204__));
  buf1  g1673(.din(new_new_n861__), .dout(new_new_n2205__));
  buf1  g1674(.din(new_new_n2205__), .dout(new_new_n2206__));
  buf1  g1675(.din(new_new_n863__), .dout(new_new_n2207__));
  buf1  g1676(.din(new_new_n2207__), .dout(new_new_n2208__));
  buf1  g1677(.din(new_new_n860__), .dout(new_new_n2209__));
  buf1  g1678(.din(new_new_n866__), .dout(new_new_n2210__));
  buf1  g1679(.din(new_new_n865__), .dout(new_new_n2211__));
  buf1  g1680(.din(new_new_n2211__), .dout(new_new_n2212__));
  buf1  g1681(.din(new_new_n867__), .dout(new_new_n2213__));
  buf1  g1682(.din(new_new_n2213__), .dout(new_new_n2214__));
  buf1  g1683(.din(new_new_n864__), .dout(new_new_n2215__));
  buf1  g1684(.din(new_new_n870__), .dout(new_new_n2216__));
  buf1  g1685(.din(new_new_n869__), .dout(new_new_n2217__));
  buf1  g1686(.din(new_new_n2217__), .dout(new_new_n2218__));
  buf1  g1687(.din(new_new_n871__), .dout(new_new_n2219__));
  buf1  g1688(.din(new_new_n2219__), .dout(new_new_n2220__));
  buf1  g1689(.din(new_new_n868__), .dout(new_new_n2221__));
  buf1  g1690(.din(new_new_n874__), .dout(new_new_n2222__));
  buf1  g1691(.din(new_new_n873__), .dout(new_new_n2223__));
  buf1  g1692(.din(new_new_n2223__), .dout(new_new_n2224__));
  buf1  g1693(.din(new_new_n875__), .dout(new_new_n2225__));
  buf1  g1694(.din(new_new_n2225__), .dout(new_new_n2226__));
  buf1  g1695(.din(new_new_n872__), .dout(new_new_n2227__));
  buf1  g1696(.din(new_new_n878__), .dout(new_new_n2228__));
  buf1  g1697(.din(new_new_n877__), .dout(new_new_n2229__));
  buf1  g1698(.din(new_new_n2229__), .dout(new_new_n2230__));
  buf1  g1699(.din(new_new_n879__), .dout(new_new_n2231__));
  buf1  g1700(.din(new_new_n2231__), .dout(new_new_n2232__));
  buf1  g1701(.din(new_new_n876__), .dout(new_new_n2233__));
  buf1  g1702(.din(new_new_n882__), .dout(new_new_n2234__));
  buf1  g1703(.din(new_new_n881__), .dout(new_new_n2235__));
  buf1  g1704(.din(new_new_n2235__), .dout(new_new_n2236__));
  buf1  g1705(.din(new_new_n883__), .dout(new_new_n2237__));
  buf1  g1706(.din(new_new_n2237__), .dout(new_new_n2238__));
  buf1  g1707(.din(new_new_n880__), .dout(new_new_n2239__));
  buf1  g1708(.din(new_new_n886__), .dout(new_new_n2240__));
  buf1  g1709(.din(new_new_n885__), .dout(new_new_n2241__));
  buf1  g1710(.din(new_new_n2241__), .dout(new_new_n2242__));
  buf1  g1711(.din(new_new_n887__), .dout(new_new_n2243__));
  buf1  g1712(.din(new_new_n2243__), .dout(new_new_n2244__));
  buf1  g1713(.din(new_new_n884__), .dout(new_new_n2245__));
  buf1  g1714(.din(new_new_n890__), .dout(new_new_n2246__));
  buf1  g1715(.din(new_new_n889__), .dout(new_new_n2247__));
  buf1  g1716(.din(new_new_n2247__), .dout(new_new_n2248__));
  buf1  g1717(.din(new_new_n891__), .dout(new_new_n2249__));
  buf1  g1718(.din(new_new_n2249__), .dout(new_new_n2250__));
  buf1  g1719(.din(new_new_n888__), .dout(new_new_n2251__));
  buf1  g1720(.din(new_new_n894__), .dout(new_new_n2252__));
  buf1  g1721(.din(new_new_n893__), .dout(new_new_n2253__));
  buf1  g1722(.din(new_new_n2253__), .dout(new_new_n2254__));
  buf1  g1723(.din(new_new_n895__), .dout(new_new_n2255__));
  buf1  g1724(.din(new_new_n2255__), .dout(new_new_n2256__));
  buf1  g1725(.din(new_new_n892__), .dout(new_new_n2257__));
  buf1  g1726(.din(new_new_n898__), .dout(new_new_n2258__));
  buf1  g1727(.din(new_new_n897__), .dout(new_new_n2259__));
  buf1  g1728(.din(new_new_n2259__), .dout(new_new_n2260__));
  buf1  g1729(.din(new_new_n899__), .dout(new_new_n2261__));
  buf1  g1730(.din(new_new_n2261__), .dout(new_new_n2262__));
  buf1  g1731(.din(new_new_n896__), .dout(new_new_n2263__));
  buf1  g1732(.din(new_new_n902__), .dout(new_new_n2264__));
  buf1  g1733(.din(new_new_n901__), .dout(new_new_n2265__));
  buf1  g1734(.din(new_new_n2265__), .dout(new_new_n2266__));
  buf1  g1735(.din(new_new_n903__), .dout(new_new_n2267__));
  buf1  g1736(.din(new_new_n2267__), .dout(new_new_n2268__));
  buf1  g1737(.din(new_new_n900__), .dout(new_new_n2269__));
  buf1  g1738(.din(new_new_n906__), .dout(new_new_n2270__));
  buf1  g1739(.din(new_new_n905__), .dout(new_new_n2271__));
  buf1  g1740(.din(new_new_n2271__), .dout(new_new_n2272__));
  buf1  g1741(.din(new_new_n907__), .dout(new_new_n2273__));
  buf1  g1742(.din(new_new_n2273__), .dout(new_new_n2274__));
  buf1  g1743(.din(new_new_n904__), .dout(new_new_n2275__));
  always @ (posedge clock) begin
    n286_lo <= n3791;
    n298_lo <= n3794;
    n310_lo <= n3797;
    n322_lo <= n3800;
    n334_lo <= n3803;
    n346_lo <= n3806;
    n358_lo <= n3809;
    n370_lo <= n3812;
    n382_lo <= n3815;
    n394_lo <= n3818;
    n406_lo <= n3821;
    n418_lo <= n3824;
    n430_lo <= n3827;
    n442_lo <= n3830;
    n454_lo <= n3833;
    n466_lo <= n3836;
    n478_lo <= n3839;
    n490_lo <= n3842;
    n502_lo <= n3845;
    n514_lo <= n3848;
    n526_lo <= n3851;
    n538_lo <= n3854;
    n550_lo <= n3857;
    n562_lo <= n3860;
    n574_lo <= n3863;
    n586_lo <= n3866;
    n598_lo <= n3869;
    n610_lo <= n3872;
    n622_lo <= n3875;
    n634_lo <= n3878;
    n646_lo <= n3881;
    n658_lo <= n3884;
    n661_lo <= n3887;
    n673_lo <= n3890;
    n685_lo <= n3893;
    n697_lo <= n3896;
    n709_lo <= n3899;
    n721_lo <= n3902;
    n733_lo <= n3905;
    n745_lo <= n3908;
    n757_lo <= n3911;
    n1248_o2 <= n3914;
    n1249_o2 <= n3917;
    n1250_o2 <= n3920;
    n1251_o2 <= n3923;
    n1252_o2 <= n3926;
    n1253_o2 <= n3929;
    n1254_o2 <= n3932;
    n1255_o2 <= n3935;
    n1207_o2 <= n3938;
    n1208_o2 <= n3941;
    n1209_o2 <= n3944;
    n1210_o2 <= n3947;
    n1211_o2 <= n3950;
    n1212_o2 <= n3953;
    n1213_o2 <= n3956;
    n1214_o2 <= n3959;
    n1215_o2 <= n3962;
    n1216_o2 <= n3965;
    n1217_o2 <= n3968;
    n1218_o2 <= n3971;
    n1219_o2 <= n3974;
    n1220_o2 <= n3977;
    n1221_o2 <= n3980;
    n1222_o2 <= n3983;
    n1223_o2 <= n3986;
    n1224_o2 <= n3989;
    n1225_o2 <= n3992;
    n1226_o2 <= n3995;
    n1227_o2 <= n3998;
    n1228_o2 <= n4001;
    n1229_o2 <= n4004;
    n1230_o2 <= n4007;
    n1231_o2 <= n4010;
    n1232_o2 <= n4013;
    n1233_o2 <= n4016;
    n1234_o2 <= n4019;
    n1235_o2 <= n4022;
    n1236_o2 <= n4025;
    n1237_o2 <= n4028;
    n1238_o2 <= n4031;
    G374_o2 <= n4034;
    G376_o2 <= n4037;
    G370_o2 <= n4040;
    G372_o2 <= n4043;
    G373_o2 <= n4046;
    G377_o2 <= n4049;
    G371_o2 <= n4052;
    G375_o2 <= n4055;
    G354_o2 <= n4058;
    G356_o2 <= n4061;
    G350_o2 <= n4064;
    G352_o2 <= n4067;
    G353_o2 <= n4070;
    G357_o2 <= n4073;
    G351_o2 <= n4076;
    G355_o2 <= n4079;
    G386_o2 <= n4082;
    G391_o2 <= n4085;
    n283_lo_buf_o2 <= n4088;
    n295_lo_buf_o2 <= n4091;
    n307_lo_buf_o2 <= n4094;
    n319_lo_buf_o2 <= n4097;
    n331_lo_buf_o2 <= n4100;
    n343_lo_buf_o2 <= n4103;
    n355_lo_buf_o2 <= n4106;
    n367_lo_buf_o2 <= n4109;
    n379_lo_buf_o2 <= n4112;
    n391_lo_buf_o2 <= n4115;
    n403_lo_buf_o2 <= n4118;
    n415_lo_buf_o2 <= n4121;
    n427_lo_buf_o2 <= n4124;
    n439_lo_buf_o2 <= n4127;
    n451_lo_buf_o2 <= n4130;
    n463_lo_buf_o2 <= n4133;
    n475_lo_buf_o2 <= n4136;
    n487_lo_buf_o2 <= n4139;
    n499_lo_buf_o2 <= n4142;
    n511_lo_buf_o2 <= n4145;
    n523_lo_buf_o2 <= n4148;
    n535_lo_buf_o2 <= n4151;
    n547_lo_buf_o2 <= n4154;
    n559_lo_buf_o2 <= n4157;
    n571_lo_buf_o2 <= n4160;
    n583_lo_buf_o2 <= n4163;
    n595_lo_buf_o2 <= n4166;
    n607_lo_buf_o2 <= n4169;
    n619_lo_buf_o2 <= n4172;
    n631_lo_buf_o2 <= n4175;
    n643_lo_buf_o2 <= n4178;
    n655_lo_buf_o2 <= n4181;
    G234_o2 <= n4184;
    G247_o2 <= n4187;
    G260_o2 <= n4190;
    G273_o2 <= n4193;
    G286_o2 <= n4196;
    G299_o2 <= n4199;
    G312_o2 <= n4202;
    G325_o2 <= n4205;
    n667_lo_buf_o2 <= n4208;
    n679_lo_buf_o2 <= n4211;
    n691_lo_buf_o2 <= n4214;
    n703_lo_buf_o2 <= n4217;
    n715_lo_buf_o2 <= n4220;
    n727_lo_buf_o2 <= n4223;
    n739_lo_buf_o2 <= n4226;
    n751_lo_buf_o2 <= n4229;
    n763_lo_buf_o2 <= n4232;
    G186_o2 <= n4235;
    G189_o2 <= n4238;
    G192_o2 <= n4241;
    G195_o2 <= n4244;
    G198_o2 <= n4247;
    G201_o2 <= n4250;
    G204_o2 <= n4253;
    G207_o2 <= n4256;
    n280_lo_buf_o2 <= n4259;
    n292_lo_buf_o2 <= n4262;
    n304_lo_buf_o2 <= n4265;
    n316_lo_buf_o2 <= n4268;
    n328_lo_buf_o2 <= n4271;
    n340_lo_buf_o2 <= n4274;
    n352_lo_buf_o2 <= n4277;
    n364_lo_buf_o2 <= n4280;
    n376_lo_buf_o2 <= n4283;
    n388_lo_buf_o2 <= n4286;
    n400_lo_buf_o2 <= n4289;
    n412_lo_buf_o2 <= n4292;
    n424_lo_buf_o2 <= n4295;
    n436_lo_buf_o2 <= n4298;
    n448_lo_buf_o2 <= n4301;
    n460_lo_buf_o2 <= n4304;
    n472_lo_buf_o2 <= n4307;
    n484_lo_buf_o2 <= n4310;
    n496_lo_buf_o2 <= n4313;
    n508_lo_buf_o2 <= n4316;
    n520_lo_buf_o2 <= n4319;
    n532_lo_buf_o2 <= n4322;
    n544_lo_buf_o2 <= n4325;
    n556_lo_buf_o2 <= n4328;
    n568_lo_buf_o2 <= n4331;
    n580_lo_buf_o2 <= n4334;
    n592_lo_buf_o2 <= n4337;
    n604_lo_buf_o2 <= n4340;
    n616_lo_buf_o2 <= n4343;
    n628_lo_buf_o2 <= n4346;
    n640_lo_buf_o2 <= n4349;
    n652_lo_buf_o2 <= n4352;
  end
  initial begin
    n286_lo <= 1'b0;
    n298_lo <= 1'b0;
    n310_lo <= 1'b0;
    n322_lo <= 1'b0;
    n334_lo <= 1'b0;
    n346_lo <= 1'b0;
    n358_lo <= 1'b0;
    n370_lo <= 1'b0;
    n382_lo <= 1'b0;
    n394_lo <= 1'b0;
    n406_lo <= 1'b0;
    n418_lo <= 1'b0;
    n430_lo <= 1'b0;
    n442_lo <= 1'b0;
    n454_lo <= 1'b0;
    n466_lo <= 1'b0;
    n478_lo <= 1'b0;
    n490_lo <= 1'b0;
    n502_lo <= 1'b0;
    n514_lo <= 1'b0;
    n526_lo <= 1'b0;
    n538_lo <= 1'b0;
    n550_lo <= 1'b0;
    n562_lo <= 1'b0;
    n574_lo <= 1'b0;
    n586_lo <= 1'b0;
    n598_lo <= 1'b0;
    n610_lo <= 1'b0;
    n622_lo <= 1'b0;
    n634_lo <= 1'b0;
    n646_lo <= 1'b0;
    n658_lo <= 1'b0;
    n661_lo <= 1'b0;
    n673_lo <= 1'b0;
    n685_lo <= 1'b0;
    n697_lo <= 1'b0;
    n709_lo <= 1'b0;
    n721_lo <= 1'b0;
    n733_lo <= 1'b0;
    n745_lo <= 1'b0;
    n757_lo <= 1'b0;
    n1248_o2 <= 1'b0;
    n1249_o2 <= 1'b0;
    n1250_o2 <= 1'b0;
    n1251_o2 <= 1'b0;
    n1252_o2 <= 1'b0;
    n1253_o2 <= 1'b0;
    n1254_o2 <= 1'b0;
    n1255_o2 <= 1'b0;
    n1207_o2 <= 1'b0;
    n1208_o2 <= 1'b0;
    n1209_o2 <= 1'b0;
    n1210_o2 <= 1'b0;
    n1211_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1213_o2 <= 1'b0;
    n1214_o2 <= 1'b0;
    n1215_o2 <= 1'b0;
    n1216_o2 <= 1'b0;
    n1217_o2 <= 1'b0;
    n1218_o2 <= 1'b0;
    n1219_o2 <= 1'b0;
    n1220_o2 <= 1'b0;
    n1221_o2 <= 1'b0;
    n1222_o2 <= 1'b0;
    n1223_o2 <= 1'b0;
    n1224_o2 <= 1'b0;
    n1225_o2 <= 1'b0;
    n1226_o2 <= 1'b0;
    n1227_o2 <= 1'b0;
    n1228_o2 <= 1'b0;
    n1229_o2 <= 1'b0;
    n1230_o2 <= 1'b0;
    n1231_o2 <= 1'b0;
    n1232_o2 <= 1'b0;
    n1233_o2 <= 1'b0;
    n1234_o2 <= 1'b0;
    n1235_o2 <= 1'b0;
    n1236_o2 <= 1'b0;
    n1237_o2 <= 1'b0;
    n1238_o2 <= 1'b0;
    G374_o2 <= 1'b0;
    G376_o2 <= 1'b0;
    G370_o2 <= 1'b0;
    G372_o2 <= 1'b0;
    G373_o2 <= 1'b0;
    G377_o2 <= 1'b0;
    G371_o2 <= 1'b0;
    G375_o2 <= 1'b0;
    G354_o2 <= 1'b0;
    G356_o2 <= 1'b0;
    G350_o2 <= 1'b0;
    G352_o2 <= 1'b0;
    G353_o2 <= 1'b0;
    G357_o2 <= 1'b0;
    G351_o2 <= 1'b0;
    G355_o2 <= 1'b0;
    G386_o2 <= 1'b0;
    G391_o2 <= 1'b0;
    n283_lo_buf_o2 <= 1'b0;
    n295_lo_buf_o2 <= 1'b0;
    n307_lo_buf_o2 <= 1'b0;
    n319_lo_buf_o2 <= 1'b0;
    n331_lo_buf_o2 <= 1'b0;
    n343_lo_buf_o2 <= 1'b0;
    n355_lo_buf_o2 <= 1'b0;
    n367_lo_buf_o2 <= 1'b0;
    n379_lo_buf_o2 <= 1'b0;
    n391_lo_buf_o2 <= 1'b0;
    n403_lo_buf_o2 <= 1'b0;
    n415_lo_buf_o2 <= 1'b0;
    n427_lo_buf_o2 <= 1'b0;
    n439_lo_buf_o2 <= 1'b0;
    n451_lo_buf_o2 <= 1'b0;
    n463_lo_buf_o2 <= 1'b0;
    n475_lo_buf_o2 <= 1'b0;
    n487_lo_buf_o2 <= 1'b0;
    n499_lo_buf_o2 <= 1'b0;
    n511_lo_buf_o2 <= 1'b0;
    n523_lo_buf_o2 <= 1'b0;
    n535_lo_buf_o2 <= 1'b0;
    n547_lo_buf_o2 <= 1'b0;
    n559_lo_buf_o2 <= 1'b0;
    n571_lo_buf_o2 <= 1'b0;
    n583_lo_buf_o2 <= 1'b0;
    n595_lo_buf_o2 <= 1'b0;
    n607_lo_buf_o2 <= 1'b0;
    n619_lo_buf_o2 <= 1'b0;
    n631_lo_buf_o2 <= 1'b0;
    n643_lo_buf_o2 <= 1'b0;
    n655_lo_buf_o2 <= 1'b0;
    G234_o2 <= 1'b0;
    G247_o2 <= 1'b0;
    G260_o2 <= 1'b0;
    G273_o2 <= 1'b0;
    G286_o2 <= 1'b0;
    G299_o2 <= 1'b0;
    G312_o2 <= 1'b0;
    G325_o2 <= 1'b0;
    n667_lo_buf_o2 <= 1'b0;
    n679_lo_buf_o2 <= 1'b0;
    n691_lo_buf_o2 <= 1'b0;
    n703_lo_buf_o2 <= 1'b0;
    n715_lo_buf_o2 <= 1'b0;
    n727_lo_buf_o2 <= 1'b0;
    n739_lo_buf_o2 <= 1'b0;
    n751_lo_buf_o2 <= 1'b0;
    n763_lo_buf_o2 <= 1'b0;
    G186_o2 <= 1'b0;
    G189_o2 <= 1'b0;
    G192_o2 <= 1'b0;
    G195_o2 <= 1'b0;
    G198_o2 <= 1'b0;
    G201_o2 <= 1'b0;
    G204_o2 <= 1'b0;
    G207_o2 <= 1'b0;
    n280_lo_buf_o2 <= 1'b0;
    n292_lo_buf_o2 <= 1'b0;
    n304_lo_buf_o2 <= 1'b0;
    n316_lo_buf_o2 <= 1'b0;
    n328_lo_buf_o2 <= 1'b0;
    n340_lo_buf_o2 <= 1'b0;
    n352_lo_buf_o2 <= 1'b0;
    n364_lo_buf_o2 <= 1'b0;
    n376_lo_buf_o2 <= 1'b0;
    n388_lo_buf_o2 <= 1'b0;
    n400_lo_buf_o2 <= 1'b0;
    n412_lo_buf_o2 <= 1'b0;
    n424_lo_buf_o2 <= 1'b0;
    n436_lo_buf_o2 <= 1'b0;
    n448_lo_buf_o2 <= 1'b0;
    n460_lo_buf_o2 <= 1'b0;
    n472_lo_buf_o2 <= 1'b0;
    n484_lo_buf_o2 <= 1'b0;
    n496_lo_buf_o2 <= 1'b0;
    n508_lo_buf_o2 <= 1'b0;
    n520_lo_buf_o2 <= 1'b0;
    n532_lo_buf_o2 <= 1'b0;
    n544_lo_buf_o2 <= 1'b0;
    n556_lo_buf_o2 <= 1'b0;
    n568_lo_buf_o2 <= 1'b0;
    n580_lo_buf_o2 <= 1'b0;
    n592_lo_buf_o2 <= 1'b0;
    n604_lo_buf_o2 <= 1'b0;
    n616_lo_buf_o2 <= 1'b0;
    n628_lo_buf_o2 <= 1'b0;
    n640_lo_buf_o2 <= 1'b0;
    n652_lo_buf_o2 <= 1'b0;
  end
endmodule


