
module mymod
(
  a_0_,
  a_1_,
  a_2_,
  a_3_,
  a_4_,
  a_5_,
  a_6_,
  a_7_,
  b_0_,
  b_1_,
  b_2_,
  b_3_,
  b_4_,
  b_5_,
  b_6_,
  b_7_,
  product_0_,
  product_1_,
  product_2_,
  product_3_,
  product_4_,
  product_5_,
  product_6_,
  product_7_
);

  input a_0_;input a_1_;input a_2_;input a_3_;input a_4_;input a_5_;input a_6_;input a_7_;input b_0_;input b_1_;input b_2_;input b_3_;input b_4_;input b_5_;input b_6_;input b_7_;
  output product_0_;output product_1_;output product_2_;output product_3_;output product_4_;output product_5_;output product_6_;output product_7_;
  wire a_0__p;
  wire a_0__n;
  wire a_1__p;
  wire a_1__n;
  wire a_2__p;
  wire a_2__n;
  wire a_3__p;
  wire a_3__n;
  wire a_4__p;
  wire a_4__n;
  wire a_5__p;
  wire a_5__n;
  wire a_6__p;
  wire a_6__n;
  wire a_7__p;
  wire a_7__n;
  wire b_0__p;
  wire b_0__n;
  wire b_1__p;
  wire b_1__n;
  wire b_2__p;
  wire b_2__n;
  wire b_3__p;
  wire b_3__n;
  wire b_4__p;
  wire b_4__n;
  wire b_5__p;
  wire b_5__n;
  wire b_6__p;
  wire b_6__n;
  wire b_7__p;
  wire b_7__n;
  wire g17_p;
  wire g17_n;
  wire g18_p;
  wire g18_n;
  wire g19_p;
  wire g19_n;
  wire g20_p;
  wire g20_n;
  wire g21_p;
  wire g21_n;
  wire g22_p;
  wire g22_n;
  wire g23_p;
  wire g23_n;
  wire g24_p;
  wire g24_n;
  wire g25_p;
  wire g25_n;
  wire g26_p;
  wire g26_n;
  wire g27_p;
  wire g27_n;
  wire g28_p;
  wire g28_n;
  wire g29_p;
  wire g29_n;
  wire g30_p;
  wire g30_n;
  wire g31_p;
  wire g31_n;
  wire g32_p;
  wire g32_n;
  wire g33_p;
  wire g33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire a_7__p_spl_;
  wire a_7__p_spl_0;
  wire a_7__p_spl_00;
  wire a_7__p_spl_01;
  wire a_7__p_spl_1;
  wire a_7__p_spl_10;
  wire a_7__p_spl_11;
  wire b_4__p_spl_;
  wire b_4__p_spl_0;
  wire b_4__p_spl_00;
  wire b_4__p_spl_01;
  wire b_4__p_spl_1;
  wire b_4__p_spl_10;
  wire b_4__p_spl_11;
  wire a_7__n_spl_;
  wire a_7__n_spl_0;
  wire a_7__n_spl_00;
  wire a_7__n_spl_01;
  wire a_7__n_spl_1;
  wire a_7__n_spl_10;
  wire a_7__n_spl_11;
  wire b_4__n_spl_;
  wire b_4__n_spl_0;
  wire b_4__n_spl_00;
  wire b_4__n_spl_01;
  wire b_4__n_spl_1;
  wire b_4__n_spl_10;
  wire b_4__n_spl_11;
  wire b_3__p_spl_;
  wire b_3__p_spl_0;
  wire b_3__p_spl_00;
  wire b_3__p_spl_000;
  wire b_3__p_spl_01;
  wire b_3__p_spl_1;
  wire b_3__p_spl_10;
  wire b_3__p_spl_11;
  wire g17_p_spl_;
  wire g17_p_spl_0;
  wire b_3__n_spl_;
  wire b_3__n_spl_0;
  wire b_3__n_spl_00;
  wire b_3__n_spl_000;
  wire b_3__n_spl_01;
  wire b_3__n_spl_1;
  wire b_3__n_spl_10;
  wire b_3__n_spl_11;
  wire g17_n_spl_;
  wire g17_n_spl_0;
  wire g19_n_spl_;
  wire g19_p_spl_;
  wire g18_n_spl_;
  wire g18_n_spl_0;
  wire g18_p_spl_;
  wire g18_p_spl_0;
  wire b_5__p_spl_;
  wire b_5__p_spl_0;
  wire b_5__p_spl_00;
  wire b_5__p_spl_01;
  wire b_5__p_spl_1;
  wire b_5__p_spl_10;
  wire b_5__p_spl_11;
  wire b_5__n_spl_;
  wire b_5__n_spl_0;
  wire b_5__n_spl_00;
  wire b_5__n_spl_01;
  wire b_5__n_spl_1;
  wire b_5__n_spl_10;
  wire b_5__n_spl_11;
  wire g21_p_spl_;
  wire g21_p_spl_0;
  wire g21_p_spl_1;
  wire g22_p_spl_;
  wire g21_n_spl_;
  wire g21_n_spl_0;
  wire g21_n_spl_1;
  wire g22_n_spl_;
  wire g23_n_spl_;
  wire g23_p_spl_;
  wire b_6__p_spl_;
  wire b_6__p_spl_0;
  wire b_6__p_spl_00;
  wire b_6__p_spl_01;
  wire b_6__p_spl_1;
  wire b_6__p_spl_10;
  wire b_6__p_spl_11;
  wire b_6__n_spl_;
  wire b_6__n_spl_0;
  wire b_6__n_spl_00;
  wire b_6__n_spl_01;
  wire b_6__n_spl_1;
  wire b_6__n_spl_10;
  wire b_6__n_spl_11;
  wire a_6__n_spl_;
  wire a_6__n_spl_0;
  wire a_6__n_spl_00;
  wire a_6__n_spl_01;
  wire a_6__n_spl_1;
  wire a_6__n_spl_10;
  wire a_6__n_spl_11;
  wire b_7__p_spl_;
  wire b_7__p_spl_0;
  wire b_7__p_spl_00;
  wire b_7__p_spl_000;
  wire b_7__p_spl_001;
  wire b_7__p_spl_01;
  wire b_7__p_spl_1;
  wire b_7__p_spl_10;
  wire b_7__p_spl_11;
  wire a_6__p_spl_;
  wire a_6__p_spl_0;
  wire a_6__p_spl_00;
  wire a_6__p_spl_01;
  wire a_6__p_spl_1;
  wire a_6__p_spl_10;
  wire a_6__p_spl_11;
  wire b_7__n_spl_;
  wire b_7__n_spl_0;
  wire b_7__n_spl_00;
  wire b_7__n_spl_000;
  wire b_7__n_spl_001;
  wire b_7__n_spl_01;
  wire b_7__n_spl_1;
  wire b_7__n_spl_10;
  wire b_7__n_spl_11;
  wire g25_p_spl_;
  wire g26_n_spl_;
  wire g25_n_spl_;
  wire g26_p_spl_;
  wire g27_n_spl_;
  wire g27_p_spl_;
  wire g24_p_spl_;
  wire g24_p_spl_0;
  wire g24_p_spl_1;
  wire g29_p_spl_;
  wire g24_n_spl_;
  wire g24_n_spl_0;
  wire g24_n_spl_1;
  wire g29_n_spl_;
  wire b_0__p_spl_;
  wire b_0__p_spl_0;
  wire b_0__p_spl_00;
  wire b_0__p_spl_000;
  wire b_0__p_spl_01;
  wire b_0__p_spl_1;
  wire b_0__p_spl_10;
  wire b_0__p_spl_11;
  wire b_0__n_spl_;
  wire b_0__n_spl_0;
  wire b_0__n_spl_00;
  wire b_0__n_spl_01;
  wire b_0__n_spl_1;
  wire b_0__n_spl_10;
  wire b_0__n_spl_11;
  wire b_1__p_spl_;
  wire b_1__p_spl_0;
  wire b_1__p_spl_00;
  wire b_1__p_spl_000;
  wire b_1__p_spl_01;
  wire b_1__p_spl_1;
  wire b_1__p_spl_10;
  wire b_1__p_spl_11;
  wire g33_p_spl_;
  wire g33_p_spl_0;
  wire b_1__n_spl_;
  wire b_1__n_spl_0;
  wire b_1__n_spl_00;
  wire b_1__n_spl_01;
  wire b_1__n_spl_1;
  wire b_1__n_spl_10;
  wire b_1__n_spl_11;
  wire g33_n_spl_;
  wire g33_n_spl_0;
  wire b_2__p_spl_;
  wire b_2__p_spl_0;
  wire b_2__p_spl_00;
  wire b_2__p_spl_000;
  wire b_2__p_spl_01;
  wire b_2__p_spl_1;
  wire b_2__p_spl_10;
  wire b_2__p_spl_11;
  wire g34_p_spl_;
  wire g34_p_spl_0;
  wire b_2__n_spl_;
  wire b_2__n_spl_0;
  wire b_2__n_spl_00;
  wire b_2__n_spl_000;
  wire b_2__n_spl_01;
  wire b_2__n_spl_1;
  wire b_2__n_spl_10;
  wire b_2__n_spl_11;
  wire g34_n_spl_;
  wire g34_n_spl_0;
  wire g32_p_spl_;
  wire g32_p_spl_0;
  wire g35_p_spl_;
  wire g35_p_spl_0;
  wire g35_p_spl_00;
  wire g35_p_spl_01;
  wire g35_p_spl_1;
  wire g35_p_spl_10;
  wire g32_n_spl_;
  wire g32_n_spl_0;
  wire g35_n_spl_;
  wire g35_n_spl_0;
  wire g35_n_spl_00;
  wire g35_n_spl_01;
  wire g35_n_spl_1;
  wire g35_n_spl_10;
  wire g37_n_spl_;
  wire g39_n_spl_;
  wire g39_n_spl_0;
  wire g37_p_spl_;
  wire g39_p_spl_;
  wire g39_p_spl_0;
  wire g40_n_spl_;
  wire g40_p_spl_;
  wire g41_n_spl_;
  wire g41_n_spl_0;
  wire g41_n_spl_00;
  wire g41_n_spl_01;
  wire g41_n_spl_1;
  wire g41_p_spl_;
  wire g41_p_spl_0;
  wire g41_p_spl_00;
  wire g41_p_spl_01;
  wire g41_p_spl_1;
  wire g42_p_spl_;
  wire g42_n_spl_;
  wire g36_n_spl_;
  wire g36_n_spl_0;
  wire g36_p_spl_;
  wire g30_p_spl_;
  wire g30_p_spl_0;
  wire g44_p_spl_;
  wire g44_p_spl_0;
  wire g44_p_spl_1;
  wire g46_n_spl_;
  wire g44_n_spl_;
  wire g44_n_spl_0;
  wire g44_n_spl_1;
  wire g46_p_spl_;
  wire g47_n_spl_;
  wire g48_p_spl_;
  wire g52_p_spl_;
  wire g52_n_spl_;
  wire g53_n_spl_;
  wire g53_p_spl_;
  wire g55_p_spl_;
  wire g55_n_spl_;
  wire g56_n_spl_;
  wire g56_p_spl_;
  wire g51_p_spl_;
  wire g57_n_spl_;
  wire g51_n_spl_;
  wire g57_p_spl_;
  wire a_5__p_spl_;
  wire a_5__p_spl_0;
  wire a_5__p_spl_00;
  wire a_5__p_spl_01;
  wire a_5__p_spl_1;
  wire a_5__p_spl_10;
  wire a_5__p_spl_11;
  wire a_5__n_spl_;
  wire a_5__n_spl_0;
  wire a_5__n_spl_00;
  wire a_5__n_spl_01;
  wire a_5__n_spl_1;
  wire a_5__n_spl_10;
  wire a_5__n_spl_11;
  wire a_4__n_spl_;
  wire a_4__n_spl_0;
  wire a_4__n_spl_00;
  wire a_4__n_spl_01;
  wire a_4__n_spl_1;
  wire a_4__n_spl_10;
  wire a_4__n_spl_11;
  wire a_4__p_spl_;
  wire a_4__p_spl_0;
  wire a_4__p_spl_00;
  wire a_4__p_spl_01;
  wire a_4__p_spl_1;
  wire a_4__p_spl_10;
  wire a_4__p_spl_11;
  wire g59_p_spl_;
  wire g60_p_spl_;
  wire g59_n_spl_;
  wire g60_n_spl_;
  wire g63_p_spl_;
  wire g64_p_spl_;
  wire g63_n_spl_;
  wire g64_n_spl_;
  wire g65_n_spl_;
  wire g65_n_spl_0;
  wire g65_p_spl_;
  wire g65_p_spl_0;
  wire g62_n_spl_;
  wire g67_p_spl_;
  wire g62_p_spl_;
  wire g67_n_spl_;
  wire g68_n_spl_;
  wire g68_p_spl_;
  wire g61_p_spl_;
  wire g61_p_spl_0;
  wire g70_p_spl_;
  wire g61_n_spl_;
  wire g61_n_spl_0;
  wire g70_n_spl_;
  wire g71_n_spl_;
  wire g71_p_spl_;
  wire g58_n_spl_;
  wire g58_p_spl_;
  wire g73_p_spl_;
  wire g75_p_spl_;
  wire g73_n_spl_;
  wire g75_n_spl_;
  wire g76_n_spl_;
  wire g76_p_spl_;
  wire g79_n_spl_;
  wire g79_p_spl_;
  wire g80_n_spl_;
  wire g80_p_spl_;
  wire g82_p_spl_;
  wire g82_n_spl_;
  wire g83_n_spl_;
  wire g83_p_spl_;
  wire g85_p_spl_;
  wire g85_n_spl_;
  wire g86_n_spl_;
  wire g86_p_spl_;
  wire g77_n_spl_;
  wire g88_p_spl_;
  wire g77_p_spl_;
  wire g88_n_spl_;
  wire g89_n_spl_;
  wire g89_p_spl_;
  wire g90_n_spl_;
  wire g92_p_spl_;
  wire g90_p_spl_;
  wire g92_n_spl_;
  wire g93_n_spl_;
  wire g93_p_spl_;
  wire g97_n_spl_;
  wire g98_n_spl_;
  wire g97_p_spl_;
  wire g98_p_spl_;
  wire g99_p_spl_;
  wire g95_n_spl_;
  wire g101_p_spl_;
  wire g95_p_spl_;
  wire g101_n_spl_;
  wire g102_p_spl_;
  wire g94_n_spl_;
  wire g104_p_spl_;
  wire g94_p_spl_;
  wire g104_n_spl_;
  wire g105_p_spl_;
  wire g109_p_spl_;
  wire g109_n_spl_;
  wire g111_n_spl_;
  wire g111_p_spl_;
  wire g110_n_spl_;
  wire g110_p_spl_;
  wire g108_p_spl_;
  wire g113_p_spl_;
  wire g108_n_spl_;
  wire g113_n_spl_;
  wire g114_n_spl_;
  wire g114_p_spl_;
  wire g116_p_spl_;
  wire g116_n_spl_;
  wire g117_n_spl_;
  wire g117_p_spl_;
  wire g118_n_spl_;
  wire g120_p_spl_;
  wire g118_p_spl_;
  wire g120_n_spl_;
  wire a_3__n_spl_;
  wire a_3__n_spl_0;
  wire a_3__n_spl_00;
  wire a_3__n_spl_01;
  wire a_3__n_spl_1;
  wire a_3__n_spl_10;
  wire a_3__n_spl_11;
  wire a_3__p_spl_;
  wire a_3__p_spl_0;
  wire a_3__p_spl_00;
  wire a_3__p_spl_01;
  wire a_3__p_spl_1;
  wire a_3__p_spl_10;
  wire a_3__p_spl_11;
  wire g122_p_spl_;
  wire g123_p_spl_;
  wire g122_n_spl_;
  wire g123_n_spl_;
  wire g125_n_spl_;
  wire g127_p_spl_;
  wire g125_p_spl_;
  wire g127_n_spl_;
  wire g128_n_spl_;
  wire g128_p_spl_;
  wire g124_p_spl_;
  wire g124_p_spl_0;
  wire g130_p_spl_;
  wire g124_n_spl_;
  wire g124_n_spl_0;
  wire g130_n_spl_;
  wire g131_n_spl_;
  wire g131_p_spl_;
  wire g121_n_spl_;
  wire g121_p_spl_;
  wire g133_p_spl_;
  wire g135_p_spl_;
  wire g133_n_spl_;
  wire g135_n_spl_;
  wire g136_n_spl_;
  wire g136_p_spl_;
  wire g137_n_spl_;
  wire g139_p_spl_;
  wire g137_p_spl_;
  wire g139_n_spl_;
  wire g140_n_spl_;
  wire g140_p_spl_;
  wire g141_n_spl_;
  wire g143_p_spl_;
  wire g141_p_spl_;
  wire g143_n_spl_;
  wire g144_n_spl_;
  wire g144_p_spl_;
  wire g145_n_spl_;
  wire g147_p_spl_;
  wire g145_p_spl_;
  wire g147_n_spl_;
  wire g151_p_spl_;
  wire g151_p_spl_0;
  wire g151_p_spl_1;
  wire g151_n_spl_;
  wire g151_n_spl_0;
  wire g151_n_spl_1;
  wire g152_n_spl_;
  wire g152_p_spl_;
  wire g150_p_spl_;
  wire g155_p_spl_;
  wire g150_n_spl_;
  wire g155_n_spl_;
  wire g156_n_spl_;
  wire g156_p_spl_;
  wire g159_n_spl_;
  wire g159_n_spl_0;
  wire g159_p_spl_;
  wire g159_p_spl_0;
  wire g158_p_spl_;
  wire g164_p_spl_;
  wire g158_n_spl_;
  wire g164_n_spl_;
  wire g165_n_spl_;
  wire g165_p_spl_;
  wire g166_n_spl_;
  wire g168_p_spl_;
  wire g166_p_spl_;
  wire g168_n_spl_;
  wire a_2__n_spl_;
  wire a_2__n_spl_0;
  wire a_2__n_spl_00;
  wire a_2__n_spl_01;
  wire a_2__n_spl_1;
  wire a_2__n_spl_10;
  wire a_2__n_spl_11;
  wire a_2__p_spl_;
  wire a_2__p_spl_0;
  wire a_2__p_spl_00;
  wire a_2__p_spl_01;
  wire a_2__p_spl_1;
  wire a_2__p_spl_10;
  wire a_2__p_spl_11;
  wire g170_p_spl_;
  wire g171_p_spl_;
  wire g170_n_spl_;
  wire g171_n_spl_;
  wire g173_n_spl_;
  wire g175_p_spl_;
  wire g173_p_spl_;
  wire g175_n_spl_;
  wire g176_n_spl_;
  wire g176_p_spl_;
  wire g172_p_spl_;
  wire g172_p_spl_0;
  wire g178_p_spl_;
  wire g172_n_spl_;
  wire g172_n_spl_0;
  wire g178_n_spl_;
  wire g179_n_spl_;
  wire g179_p_spl_;
  wire g169_n_spl_;
  wire g169_p_spl_;
  wire g181_p_spl_;
  wire g183_p_spl_;
  wire g181_n_spl_;
  wire g183_n_spl_;
  wire g184_n_spl_;
  wire g184_p_spl_;
  wire g185_n_spl_;
  wire g187_p_spl_;
  wire g185_p_spl_;
  wire g187_n_spl_;
  wire g188_n_spl_;
  wire g188_p_spl_;
  wire g189_n_spl_;
  wire g191_p_spl_;
  wire g189_p_spl_;
  wire g191_n_spl_;
  wire g192_n_spl_;
  wire g192_p_spl_;
  wire g193_n_spl_;
  wire g195_p_spl_;
  wire g193_p_spl_;
  wire g195_n_spl_;
  wire g197_n_spl_;
  wire g197_p_spl_;
  wire g198_p_spl_;
  wire g198_p_spl_0;
  wire g200_p_spl_;
  wire g198_n_spl_;
  wire g198_n_spl_0;
  wire g200_n_spl_;
  wire g201_n_spl_;
  wire g201_p_spl_;
  wire g203_p_spl_;
  wire g203_n_spl_;
  wire g202_n_spl_;
  wire g206_n_spl_;
  wire g202_p_spl_;
  wire g206_p_spl_;
  wire g209_p_spl_;
  wire g209_n_spl_;
  wire g210_n_spl_;
  wire g210_p_spl_;
  wire g208_p_spl_;
  wire g212_p_spl_;
  wire g208_n_spl_;
  wire g212_n_spl_;
  wire g213_n_spl_;
  wire g213_p_spl_;
  wire g207_n_spl_;
  wire g207_p_spl_;
  wire g215_p_spl_;
  wire g217_p_spl_;
  wire g215_n_spl_;
  wire g217_n_spl_;
  wire g218_n_spl_;
  wire g218_p_spl_;
  wire g219_n_spl_;
  wire g221_p_spl_;
  wire g219_p_spl_;
  wire g221_n_spl_;
  wire a_1__n_spl_;
  wire a_1__n_spl_0;
  wire a_1__n_spl_00;
  wire a_1__n_spl_01;
  wire a_1__n_spl_1;
  wire a_1__n_spl_10;
  wire a_1__p_spl_;
  wire a_1__p_spl_0;
  wire a_1__p_spl_00;
  wire a_1__p_spl_01;
  wire a_1__p_spl_1;
  wire a_1__p_spl_10;
  wire a_1__p_spl_11;
  wire g223_p_spl_;
  wire g223_p_spl_0;
  wire g224_p_spl_;
  wire g223_n_spl_;
  wire g223_n_spl_0;
  wire g224_n_spl_;
  wire g226_n_spl_;
  wire g228_p_spl_;
  wire g226_p_spl_;
  wire g228_n_spl_;
  wire g229_n_spl_;
  wire g229_p_spl_;
  wire g225_p_spl_;
  wire g225_p_spl_0;
  wire g231_p_spl_;
  wire g225_n_spl_;
  wire g225_n_spl_0;
  wire g231_n_spl_;
  wire g232_n_spl_;
  wire g232_p_spl_;
  wire g222_n_spl_;
  wire g222_p_spl_;
  wire g234_p_spl_;
  wire g236_p_spl_;
  wire g234_n_spl_;
  wire g236_n_spl_;
  wire g237_n_spl_;
  wire g237_p_spl_;
  wire g238_n_spl_;
  wire g240_p_spl_;
  wire g238_p_spl_;
  wire g240_n_spl_;
  wire g241_n_spl_;
  wire g241_p_spl_;
  wire g242_n_spl_;
  wire g244_p_spl_;
  wire g242_p_spl_;
  wire g244_n_spl_;
  wire g245_n_spl_;
  wire g245_p_spl_;
  wire g246_n_spl_;
  wire g248_p_spl_;
  wire g246_p_spl_;
  wire g248_n_spl_;
  wire g249_n_spl_;
  wire g249_p_spl_;
  wire g252_p_spl_;
  wire g252_p_spl_0;
  wire g252_n_spl_;
  wire g252_n_spl_0;
  wire g253_n_spl_;
  wire g253_p_spl_;
  wire g254_p_spl_;
  wire g254_p_spl_0;
  wire g258_p_spl_;
  wire g254_n_spl_;
  wire g254_n_spl_0;
  wire g258_n_spl_;
  wire g259_n_spl_;
  wire g259_p_spl_;
  wire g260_n_spl_;
  wire g262_p_spl_;
  wire g260_p_spl_;
  wire g262_n_spl_;
  wire g265_n_spl_;
  wire g265_p_spl_;
  wire g264_p_spl_;
  wire g264_p_spl_0;
  wire g269_p_spl_;
  wire g264_n_spl_;
  wire g264_n_spl_0;
  wire g269_n_spl_;
  wire g270_n_spl_;
  wire g270_p_spl_;
  wire g263_n_spl_;
  wire g263_p_spl_;
  wire g272_p_spl_;
  wire g274_p_spl_;
  wire g272_n_spl_;
  wire g274_n_spl_;
  wire g275_n_spl_;
  wire g275_p_spl_;
  wire g276_n_spl_;
  wire g278_p_spl_;
  wire g276_p_spl_;
  wire g278_n_spl_;
  wire g280_p_spl_;
  wire g280_p_spl_0;
  wire g280_n_spl_;
  wire g280_n_spl_0;
  wire a_0__n_spl_;
  wire a_0__n_spl_0;
  wire a_0__n_spl_00;
  wire a_0__n_spl_01;
  wire a_0__n_spl_1;
  wire a_0__n_spl_10;
  wire a_0__p_spl_;
  wire a_0__p_spl_0;
  wire a_0__p_spl_00;
  wire a_0__p_spl_01;
  wire a_0__p_spl_1;
  wire a_0__p_spl_10;
  wire a_0__p_spl_11;
  wire g281_n_spl_;
  wire g281_p_spl_;
  wire g282_p_spl_;
  wire g286_p_spl_;
  wire g282_n_spl_;
  wire g286_n_spl_;
  wire g287_n_spl_;
  wire g287_p_spl_;
  wire g289_n_spl_;
  wire g291_p_spl_;
  wire g289_p_spl_;
  wire g291_n_spl_;
  wire g292_n_spl_;
  wire g292_p_spl_;
  wire g288_n_spl_;
  wire g294_p_spl_;
  wire g288_p_spl_;
  wire g294_n_spl_;
  wire g295_n_spl_;
  wire g295_p_spl_;
  wire g279_n_spl_;
  wire g279_p_spl_;
  wire g297_p_spl_;
  wire g299_p_spl_;
  wire g297_n_spl_;
  wire g299_n_spl_;
  wire g300_n_spl_;
  wire g300_p_spl_;
  wire g301_n_spl_;
  wire g303_p_spl_;
  wire g301_p_spl_;
  wire g303_n_spl_;
  wire g304_n_spl_;
  wire g304_p_spl_;
  wire g305_n_spl_;
  wire g307_p_spl_;
  wire g305_p_spl_;
  wire g307_n_spl_;
  wire g308_n_spl_;
  wire g308_p_spl_;
  wire g309_n_spl_;
  wire g311_p_spl_;
  wire g309_p_spl_;
  wire g311_n_spl_;
  wire g312_n_spl_;
  wire g312_p_spl_;
  wire g315_p_spl_;
  wire g315_n_spl_;
  wire g316_n_spl_;
  wire g316_p_spl_;
  wire g317_p_spl_;
  wire g319_p_spl_;
  wire g317_n_spl_;
  wire g319_n_spl_;
  wire g320_n_spl_;
  wire g320_p_spl_;
  wire g321_n_spl_;
  wire g323_p_spl_;
  wire g321_p_spl_;
  wire g323_n_spl_;
  wire g325_p_spl_;
  wire g325_p_spl_0;
  wire g325_n_spl_;
  wire g325_n_spl_0;
  wire g326_n_spl_;
  wire g326_p_spl_;
  wire g330_p_spl_;
  wire g330_n_spl_;
  wire g331_n_spl_;
  wire g331_p_spl_;
  wire g324_n_spl_;
  wire g324_p_spl_;
  wire g333_p_spl_;
  wire g335_p_spl_;
  wire g333_n_spl_;
  wire g335_n_spl_;
  wire g336_n_spl_;
  wire g336_p_spl_;
  wire g337_n_spl_;
  wire g339_p_spl_;
  wire g337_p_spl_;
  wire g339_n_spl_;
  wire g341_n_spl_;
  wire g343_p_spl_;
  wire g341_p_spl_;
  wire g343_n_spl_;
  wire g344_n_spl_;
  wire g344_n_spl_0;
  wire g344_p_spl_;
  wire g344_p_spl_0;
  wire g340_n_spl_;
  wire g340_p_spl_;
  wire g346_p_spl_;
  wire g348_p_spl_;
  wire g346_n_spl_;
  wire g348_n_spl_;
  wire g349_n_spl_;
  wire g349_p_spl_;
  wire g350_n_spl_;
  wire g352_p_spl_;
  wire g350_p_spl_;
  wire g352_n_spl_;
  wire g353_n_spl_;
  wire g353_p_spl_;
  wire g355_p_spl_;
  wire g355_n_spl_;
  wire g356_n_spl_;
  wire g356_p_spl_;
  wire g357_n_spl_;
  wire g359_p_spl_;
  wire g357_p_spl_;
  wire g359_n_spl_;
  wire g361_p_spl_;
  wire g362_p_spl_;
  wire g362_p_spl_0;
  wire g361_n_spl_;
  wire g362_n_spl_;
  wire g362_n_spl_0;
  wire g363_n_spl_;
  wire g363_p_spl_;
  wire g364_p_spl_;
  wire g366_p_spl_;
  wire g364_n_spl_;
  wire g366_n_spl_;
  wire g367_n_spl_;
  wire g367_p_spl_;
  wire g368_n_spl_;
  wire g370_p_spl_;
  wire g368_p_spl_;
  wire g370_n_spl_;
  wire g373_p_spl_;
  wire g373_p_spl_0;
  wire g373_n_spl_;
  wire g373_n_spl_0;
  wire g374_n_spl_;
  wire g374_p_spl_;
  wire g372_p_spl_;
  wire g376_p_spl_;
  wire g372_n_spl_;
  wire g376_n_spl_;
  wire g377_n_spl_;
  wire g377_p_spl_;
  wire g371_n_spl_;
  wire g371_p_spl_;
  wire g379_p_spl_;
  wire g381_p_spl_;
  wire g379_n_spl_;
  wire g381_n_spl_;
  wire g382_n_spl_;
  wire g382_p_spl_;
  wire g383_n_spl_;
  wire g385_p_spl_;
  wire g383_p_spl_;
  wire g385_n_spl_;
  wire g387_n_spl_;
  wire g388_p_spl_;
  wire g387_p_spl_;
  wire g388_n_spl_;
  wire g389_n_spl_;
  wire g389_n_spl_0;
  wire g389_p_spl_;
  wire g389_p_spl_0;
  wire g386_n_spl_;
  wire g386_p_spl_;
  wire g391_p_spl_;
  wire g393_p_spl_;
  wire g391_n_spl_;
  wire g393_n_spl_;
  wire g394_n_spl_;
  wire g394_p_spl_;
  wire g395_n_spl_;
  wire g397_p_spl_;
  wire g395_p_spl_;
  wire g397_n_spl_;
  wire g398_n_spl_;
  wire g398_p_spl_;
  wire g400_p_spl_;
  wire g400_n_spl_;
  wire g401_n_spl_;
  wire g401_p_spl_;
  wire g402_n_spl_;
  wire g404_p_spl_;
  wire g402_p_spl_;
  wire g404_n_spl_;
  wire g406_p_spl_;
  wire g406_p_spl_0;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g407_n_spl_;
  wire g407_p_spl_;
  wire g408_p_spl_;
  wire g412_p_spl_;
  wire g408_n_spl_;
  wire g412_n_spl_;
  wire g413_n_spl_;
  wire g413_p_spl_;
  wire g414_n_spl_;
  wire g416_p_spl_;
  wire g414_p_spl_;
  wire g416_n_spl_;
  wire g418_p_spl_;
  wire g418_p_spl_0;
  wire g418_n_spl_;
  wire g418_n_spl_0;
  wire g419_n_spl_;
  wire g419_n_spl_0;
  wire g419_p_spl_;
  wire g419_p_spl_0;
  wire g417_n_spl_;
  wire g417_p_spl_;
  wire g423_p_spl_;
  wire g425_p_spl_;
  wire g423_n_spl_;
  wire g425_n_spl_;
  wire g426_n_spl_;
  wire g426_p_spl_;
  wire g427_n_spl_;
  wire g429_p_spl_;
  wire g427_p_spl_;
  wire g429_n_spl_;
  wire g430_n_spl_;
  wire g430_p_spl_;
  wire g432_p_spl_;
  wire g432_n_spl_;
  wire g433_n_spl_;
  wire g433_p_spl_;
  wire g434_n_spl_;
  wire g436_p_spl_;
  wire g434_p_spl_;
  wire g436_n_spl_;
  wire g437_p_spl_;
  wire g437_p_spl_0;
  wire g439_p_spl_;
  wire g437_n_spl_;
  wire g437_n_spl_0;
  wire g439_n_spl_;
  wire g440_n_spl_;
  wire g440_p_spl_;
  wire g445_p_spl_;
  wire g445_p_spl_0;
  wire g445_n_spl_;
  wire g445_n_spl_0;
  wire g446_n_spl_;
  wire g446_p_spl_;
  wire g447_p_spl_;
  wire g449_p_spl_;
  wire g447_n_spl_;
  wire g449_n_spl_;
  wire g450_n_spl_;
  wire g450_p_spl_;
  wire g451_n_spl_;
  wire g453_p_spl_;
  wire g451_p_spl_;
  wire g453_n_spl_;
  wire g454_n_spl_;
  wire g454_p_spl_;
  wire g456_p_spl_;
  wire g456_n_spl_;
  wire g457_n_spl_;
  wire g457_p_spl_;
  wire g458_n_spl_;
  wire g460_p_spl_;
  wire g458_p_spl_;
  wire g460_n_spl_;
  wire g461_p_spl_;
  wire g461_p_spl_0;
  wire g463_p_spl_;
  wire g463_p_spl_0;
  wire g461_n_spl_;
  wire g461_n_spl_0;
  wire g463_n_spl_;
  wire g463_n_spl_0;
  wire g465_p_spl_;
  wire g466_p_spl_;
  wire g468_p_spl_;
  wire g466_n_spl_;
  wire g469_p_spl_;
  wire g471_p_spl_;
  wire g469_n_spl_;
  wire g472_p_spl_;
  wire g474_p_spl_;
  wire g472_n_spl_;
  wire g475_p_spl_;
  wire g475_n_spl_;
  wire g475_n_spl_0;
  wire g444_p_spl_;
  wire g477_n_spl_;
  wire g442_p_spl_;
  wire g478_p_spl_;
  wire g478_n_spl_;
  wire g479_n_spl_;
  wire g405_n_spl_;
  wire g405_p_spl_;
  wire g480_n_spl_;
  wire g482_p_spl_;
  wire g483_n_spl_;
  wire g360_n_spl_;
  wire g360_p_spl_;
  wire g484_n_spl_;
  wire g486_p_spl_;
  wire g487_n_spl_;
  wire g314_p_spl_;
  wire g488_n_spl_;
  wire g489_n_spl_;
  wire g251_p_spl_;
  wire g490_n_spl_;
  wire g491_n_spl_;
  wire g196_n_spl_;
  wire g196_p_spl_;
  wire g492_n_spl_;
  wire g494_p_spl_;
  wire g495_n_spl_;
  wire g149_n_spl_;
  wire g496_n_spl_;
  wire g149_p_spl_;
  wire g496_p_spl_;
  wire g148_n_spl_;
  wire g148_p_spl_;
  wire g107_p_spl_;
  wire g498_n_spl_;
  wire g511_p_spl_;
  wire g513_p_spl_;
  wire g520_p_spl_;
  wire g522_p_spl_;
  wire g518_p_spl_;
  wire g516_p_spl_;
  wire g509_n_spl_;
  wire g505_n_spl_;
  wire g505_n_spl_0;
  wire g538_p_spl_;
  wire g538_p_spl_0;
  wire g538_p_spl_00;
  wire g538_p_spl_01;
  wire g538_p_spl_1;
  wire g538_p_spl_10;
  wire g528_n_spl_;
  wire g528_n_spl_0;
  wire g528_n_spl_00;
  wire g528_n_spl_01;
  wire g528_n_spl_1;
  wire g528_n_spl_10;

  buf

  (
    a_0__p,
    a_0_
  );


  not

  (
    a_0__n,
    a_0_
  );


  buf

  (
    a_1__p,
    a_1_
  );


  not

  (
    a_1__n,
    a_1_
  );


  buf

  (
    a_2__p,
    a_2_
  );


  not

  (
    a_2__n,
    a_2_
  );


  buf

  (
    a_3__p,
    a_3_
  );


  not

  (
    a_3__n,
    a_3_
  );


  buf

  (
    a_4__p,
    a_4_
  );


  not

  (
    a_4__n,
    a_4_
  );


  buf

  (
    a_5__p,
    a_5_
  );


  not

  (
    a_5__n,
    a_5_
  );


  buf

  (
    a_6__p,
    a_6_
  );


  not

  (
    a_6__n,
    a_6_
  );


  buf

  (
    a_7__p,
    a_7_
  );


  not

  (
    a_7__n,
    a_7_
  );


  buf

  (
    b_0__p,
    b_0_
  );


  not

  (
    b_0__n,
    b_0_
  );


  buf

  (
    b_1__p,
    b_1_
  );


  not

  (
    b_1__n,
    b_1_
  );


  buf

  (
    b_2__p,
    b_2_
  );


  not

  (
    b_2__n,
    b_2_
  );


  buf

  (
    b_3__p,
    b_3_
  );


  not

  (
    b_3__n,
    b_3_
  );


  buf

  (
    b_4__p,
    b_4_
  );


  not

  (
    b_4__n,
    b_4_
  );


  buf

  (
    b_5__p,
    b_5_
  );


  not

  (
    b_5__n,
    b_5_
  );


  buf

  (
    b_6__p,
    b_6_
  );


  not

  (
    b_6__n,
    b_6_
  );


  buf

  (
    b_7__p,
    b_7_
  );


  not

  (
    b_7__n,
    b_7_
  );


  and

  (
    g17_p,
    a_7__p_spl_00,
    b_4__p_spl_00
  );


  or

  (
    g17_n,
    a_7__n_spl_00,
    b_4__n_spl_00
  );


  and

  (
    g18_p,
    b_3__p_spl_000,
    g17_p_spl_0
  );


  or

  (
    g18_n,
    b_3__n_spl_000,
    g17_n_spl_0
  );


  and

  (
    g19_p,
    a_7__p_spl_00,
    b_3__p_spl_000
  );


  or

  (
    g19_n,
    a_7__n_spl_00,
    b_3__n_spl_000
  );


  and

  (
    g20_p,
    g17_n_spl_0,
    g19_n_spl_
  );


  or

  (
    g20_n,
    g17_p_spl_0,
    g19_p_spl_
  );


  and

  (
    g21_p,
    g18_n_spl_0,
    g20_n
  );


  or

  (
    g21_n,
    g18_p_spl_0,
    g20_p
  );


  and

  (
    g22_p,
    a_7__p_spl_01,
    b_5__p_spl_00
  );


  or

  (
    g22_n,
    a_7__n_spl_01,
    b_5__n_spl_00
  );


  and

  (
    g23_p,
    g21_p_spl_0,
    g22_p_spl_
  );


  or

  (
    g23_n,
    g21_n_spl_0,
    g22_n_spl_
  );


  and

  (
    g24_p,
    g18_n_spl_0,
    g23_n_spl_
  );


  or

  (
    g24_n,
    g18_p_spl_0,
    g23_p_spl_
  );


  and

  (
    g25_p,
    a_7__p_spl_01,
    b_6__p_spl_00
  );


  or

  (
    g25_n,
    a_7__n_spl_01,
    b_6__n_spl_00
  );


  and

  (
    g26_p,
    a_6__n_spl_00,
    b_7__p_spl_000
  );


  or

  (
    g26_n,
    a_6__p_spl_00,
    b_7__n_spl_000
  );


  and

  (
    g27_p,
    g25_p_spl_,
    g26_n_spl_
  );


  or

  (
    g27_n,
    g25_n_spl_,
    g26_p_spl_
  );


  and

  (
    g28_p,
    a_7__n_spl_10,
    b_7__p_spl_000
  );


  or

  (
    g28_n,
    a_7__p_spl_10,
    b_7__n_spl_000
  );


  and

  (
    g29_p,
    g27_n_spl_,
    g28_n
  );


  or

  (
    g29_n,
    g27_p_spl_,
    g28_p
  );


  and

  (
    g30_p,
    g24_p_spl_0,
    g29_p_spl_
  );


  or

  (
    g30_n,
    g24_n_spl_0,
    g29_n_spl_
  );


  and

  (
    g31_p,
    g21_n_spl_0,
    g22_n_spl_
  );


  or

  (
    g31_n,
    g21_p_spl_0,
    g22_p_spl_
  );


  and

  (
    g32_p,
    g23_n_spl_,
    g31_n
  );


  or

  (
    g32_n,
    g23_p_spl_,
    g31_p
  );


  and

  (
    g33_p,
    a_7__p_spl_10,
    b_0__p_spl_000
  );


  or

  (
    g33_n,
    a_7__n_spl_10,
    b_0__n_spl_00
  );


  and

  (
    g34_p,
    b_1__p_spl_000,
    g33_p_spl_0
  );


  or

  (
    g34_n,
    b_1__n_spl_00,
    g33_n_spl_0
  );


  and

  (
    g35_p,
    b_2__p_spl_000,
    g34_p_spl_0
  );


  or

  (
    g35_n,
    b_2__n_spl_000,
    g34_n_spl_0
  );


  and

  (
    g36_p,
    g32_p_spl_0,
    g35_p_spl_00
  );


  or

  (
    g36_n,
    g32_n_spl_0,
    g35_n_spl_00
  );


  and

  (
    g37_p,
    a_7__p_spl_11,
    b_2__p_spl_000
  );


  or

  (
    g37_n,
    a_7__n_spl_11,
    b_2__n_spl_000
  );


  and

  (
    g38_p,
    b_0__n_spl_00,
    b_1__n_spl_00
  );


  or

  (
    g38_n,
    b_0__p_spl_000,
    b_1__p_spl_000
  );


  and

  (
    g39_p,
    a_7__p_spl_11,
    g38_n
  );


  or

  (
    g39_n,
    a_7__n_spl_11,
    g38_p
  );


  and

  (
    g40_p,
    g37_n_spl_,
    g39_n_spl_0
  );


  or

  (
    g40_n,
    g37_p_spl_,
    g39_p_spl_0
  );


  and

  (
    g41_p,
    g35_n_spl_00,
    g40_n_spl_
  );


  or

  (
    g41_n,
    g35_p_spl_00,
    g40_p_spl_
  );


  and

  (
    g42_p,
    g32_n_spl_0,
    g41_n_spl_00
  );


  or

  (
    g42_n,
    g32_p_spl_0,
    g41_p_spl_00
  );


  and

  (
    g43_p,
    g35_n_spl_01,
    g42_p_spl_
  );


  or

  (
    g43_n,
    g35_p_spl_01,
    g42_n_spl_
  );


  and

  (
    g44_p,
    g36_n_spl_0,
    g43_n
  );


  or

  (
    g44_n,
    g36_p_spl_,
    g43_p
  );


  and

  (
    g45_p,
    g24_n_spl_0,
    g29_n_spl_
  );


  or

  (
    g45_n,
    g24_p_spl_0,
    g29_p_spl_
  );


  and

  (
    g46_p,
    g30_n,
    g45_n
  );


  or

  (
    g46_n,
    g30_p_spl_0,
    g45_p
  );


  and

  (
    g47_p,
    g44_p_spl_0,
    g46_n_spl_
  );


  or

  (
    g47_n,
    g44_n_spl_0,
    g46_p_spl_
  );


  and

  (
    g48_p,
    g36_n_spl_0,
    g47_n_spl_
  );


  and

  (
    g49_p,
    g30_p_spl_0,
    g48_p_spl_
  );


  and

  (
    g50_p,
    g32_p_spl_,
    g41_p_spl_00
  );


  or

  (
    g50_n,
    g32_n_spl_,
    g41_n_spl_00
  );


  and

  (
    g51_p,
    g42_n_spl_,
    g50_n
  );


  or

  (
    g51_n,
    g42_p_spl_,
    g50_p
  );


  and

  (
    g52_p,
    a_6__p_spl_00,
    b_5__p_spl_00
  );


  or

  (
    g52_n,
    a_6__n_spl_00,
    b_5__n_spl_00
  );


  and

  (
    g53_p,
    g21_p_spl_1,
    g52_p_spl_
  );


  or

  (
    g53_n,
    g21_n_spl_1,
    g52_n_spl_
  );


  and

  (
    g54_p,
    g21_n_spl_1,
    g52_n_spl_
  );


  or

  (
    g54_n,
    g21_p_spl_1,
    g52_p_spl_
  );


  and

  (
    g55_p,
    g53_n_spl_,
    g54_n
  );


  or

  (
    g55_n,
    g53_p_spl_,
    g54_p
  );


  and

  (
    g56_p,
    g41_p_spl_01,
    g55_p_spl_
  );


  or

  (
    g56_n,
    g41_n_spl_01,
    g55_n_spl_
  );


  and

  (
    g57_p,
    g35_n_spl_01,
    g56_n_spl_
  );


  or

  (
    g57_n,
    g35_p_spl_01,
    g56_p_spl_
  );


  and

  (
    g58_p,
    g51_p_spl_,
    g57_n_spl_
  );


  or

  (
    g58_n,
    g51_n_spl_,
    g57_p_spl_
  );


  and

  (
    g59_p,
    a_5__p_spl_00,
    b_6__p_spl_00
  );


  or

  (
    g59_n,
    a_5__n_spl_00,
    b_6__n_spl_00
  );


  and

  (
    g60_p,
    a_4__n_spl_00,
    b_7__p_spl_001
  );


  or

  (
    g60_n,
    a_4__p_spl_00,
    b_7__n_spl_001
  );


  and

  (
    g61_p,
    g59_p_spl_,
    g60_p_spl_
  );


  or

  (
    g61_n,
    g59_n_spl_,
    g60_n_spl_
  );


  and

  (
    g62_p,
    g18_n_spl_,
    g53_n_spl_
  );


  or

  (
    g62_n,
    g18_p_spl_,
    g53_p_spl_
  );


  and

  (
    g63_p,
    a_6__p_spl_01,
    b_6__p_spl_01
  );


  or

  (
    g63_n,
    a_6__n_spl_01,
    b_6__n_spl_01
  );


  and

  (
    g64_p,
    a_5__n_spl_00,
    b_7__p_spl_001
  );


  or

  (
    g64_n,
    a_5__p_spl_00,
    b_7__n_spl_001
  );


  and

  (
    g65_p,
    g63_p_spl_,
    g64_p_spl_
  );


  or

  (
    g65_n,
    g63_n_spl_,
    g64_n_spl_
  );


  and

  (
    g66_p,
    g63_n_spl_,
    g64_n_spl_
  );


  or

  (
    g66_n,
    g63_p_spl_,
    g64_p_spl_
  );


  and

  (
    g67_p,
    g65_n_spl_0,
    g66_n
  );


  or

  (
    g67_n,
    g65_p_spl_0,
    g66_p
  );


  and

  (
    g68_p,
    g62_n_spl_,
    g67_p_spl_
  );


  or

  (
    g68_n,
    g62_p_spl_,
    g67_n_spl_
  );


  and

  (
    g69_p,
    g62_p_spl_,
    g67_n_spl_
  );


  or

  (
    g69_n,
    g62_n_spl_,
    g67_p_spl_
  );


  and

  (
    g70_p,
    g68_n_spl_,
    g69_n
  );


  or

  (
    g70_n,
    g68_p_spl_,
    g69_p
  );


  and

  (
    g71_p,
    g61_p_spl_0,
    g70_p_spl_
  );


  or

  (
    g71_n,
    g61_n_spl_0,
    g70_n_spl_
  );


  and

  (
    g72_p,
    g61_n_spl_0,
    g70_n_spl_
  );


  or

  (
    g72_n,
    g61_p_spl_0,
    g70_p_spl_
  );


  and

  (
    g73_p,
    g71_n_spl_,
    g72_n
  );


  or

  (
    g73_n,
    g71_p_spl_,
    g72_p
  );


  and

  (
    g74_p,
    g51_n_spl_,
    g57_p_spl_
  );


  or

  (
    g74_n,
    g51_p_spl_,
    g57_n_spl_
  );


  and

  (
    g75_p,
    g58_n_spl_,
    g74_n
  );


  or

  (
    g75_n,
    g58_p_spl_,
    g74_p
  );


  and

  (
    g76_p,
    g73_p_spl_,
    g75_p_spl_
  );


  or

  (
    g76_n,
    g73_n_spl_,
    g75_n_spl_
  );


  and

  (
    g77_p,
    g58_n_spl_,
    g76_n_spl_
  );


  or

  (
    g77_n,
    g58_p_spl_,
    g76_p_spl_
  );


  and

  (
    g78_p,
    g25_n_spl_,
    g26_p_spl_
  );


  or

  (
    g78_n,
    g25_p_spl_,
    g26_n_spl_
  );


  and

  (
    g79_p,
    g27_n_spl_,
    g78_n
  );


  or

  (
    g79_n,
    g27_p_spl_,
    g78_p
  );


  and

  (
    g80_p,
    g24_n_spl_1,
    g79_n_spl_
  );


  or

  (
    g80_n,
    g24_p_spl_1,
    g79_p_spl_
  );


  and

  (
    g81_p,
    g24_p_spl_1,
    g79_p_spl_
  );


  or

  (
    g81_n,
    g24_n_spl_1,
    g79_n_spl_
  );


  and

  (
    g82_p,
    g80_n_spl_,
    g81_n
  );


  or

  (
    g82_n,
    g80_p_spl_,
    g81_p
  );


  and

  (
    g83_p,
    g65_p_spl_0,
    g82_p_spl_
  );


  or

  (
    g83_n,
    g65_n_spl_0,
    g82_n_spl_
  );


  and

  (
    g84_p,
    g65_n_spl_,
    g82_n_spl_
  );


  or

  (
    g84_n,
    g65_p_spl_,
    g82_p_spl_
  );


  and

  (
    g85_p,
    g83_n_spl_,
    g84_n
  );


  or

  (
    g85_n,
    g83_p_spl_,
    g84_p
  );


  and

  (
    g86_p,
    g44_p_spl_0,
    g85_p_spl_
  );


  or

  (
    g86_n,
    g44_n_spl_0,
    g85_n_spl_
  );


  and

  (
    g87_p,
    g44_n_spl_1,
    g85_n_spl_
  );


  or

  (
    g87_n,
    g44_p_spl_1,
    g85_p_spl_
  );


  and

  (
    g88_p,
    g86_n_spl_,
    g87_n
  );


  or

  (
    g88_n,
    g86_p_spl_,
    g87_p
  );


  and

  (
    g89_p,
    g77_n_spl_,
    g88_p_spl_
  );


  or

  (
    g89_n,
    g77_p_spl_,
    g88_n_spl_
  );


  and

  (
    g90_p,
    g68_n_spl_,
    g71_n_spl_
  );


  or

  (
    g90_n,
    g68_p_spl_,
    g71_p_spl_
  );


  and

  (
    g91_p,
    g77_p_spl_,
    g88_n_spl_
  );


  or

  (
    g91_n,
    g77_n_spl_,
    g88_p_spl_
  );


  and

  (
    g92_p,
    g89_n_spl_,
    g91_n
  );


  or

  (
    g92_n,
    g89_p_spl_,
    g91_p
  );


  and

  (
    g93_p,
    g90_n_spl_,
    g92_p_spl_
  );


  or

  (
    g93_n,
    g90_p_spl_,
    g92_n_spl_
  );


  and

  (
    g94_p,
    g89_n_spl_,
    g93_n_spl_
  );


  or

  (
    g94_n,
    g89_p_spl_,
    g93_p_spl_
  );


  and

  (
    g95_p,
    g80_n_spl_,
    g83_n_spl_
  );


  or

  (
    g95_n,
    g80_p_spl_,
    g83_p_spl_
  );


  and

  (
    g96_p,
    g44_n_spl_1,
    g46_p_spl_
  );


  or

  (
    g96_n,
    g44_p_spl_1,
    g46_n_spl_
  );


  and

  (
    g97_p,
    g47_n_spl_,
    g96_n
  );


  or

  (
    g97_n,
    g47_p,
    g96_p
  );


  and

  (
    g98_p,
    g36_n_spl_,
    g86_n_spl_
  );


  or

  (
    g98_n,
    g36_p_spl_,
    g86_p_spl_
  );


  and

  (
    g99_p,
    g97_n_spl_,
    g98_n_spl_
  );


  or

  (
    g99_n,
    g97_p_spl_,
    g98_p_spl_
  );


  and

  (
    g100_p,
    g97_p_spl_,
    g98_p_spl_
  );


  or

  (
    g100_n,
    g97_n_spl_,
    g98_n_spl_
  );


  and

  (
    g101_p,
    g99_n,
    g100_n
  );


  or

  (
    g101_n,
    g99_p_spl_,
    g100_p
  );


  and

  (
    g102_p,
    g95_n_spl_,
    g101_p_spl_
  );


  or

  (
    g102_n,
    g95_p_spl_,
    g101_n_spl_
  );


  and

  (
    g103_p,
    g95_p_spl_,
    g101_n_spl_
  );


  or

  (
    g103_n,
    g95_n_spl_,
    g101_p_spl_
  );


  and

  (
    g104_p,
    g102_n,
    g103_n
  );


  or

  (
    g104_n,
    g102_p_spl_,
    g103_p
  );


  and

  (
    g105_p,
    g94_n_spl_,
    g104_p_spl_
  );


  or

  (
    g105_n,
    g94_p_spl_,
    g104_n_spl_
  );


  and

  (
    g106_p,
    g94_p_spl_,
    g104_n_spl_
  );


  or

  (
    g106_n,
    g94_n_spl_,
    g104_p_spl_
  );


  and

  (
    g107_p,
    g105_n,
    g106_n
  );


  or

  (
    g107_n,
    g105_p_spl_,
    g106_p
  );


  and

  (
    g108_p,
    a_5__p_spl_01,
    b_5__p_spl_01
  );


  or

  (
    g108_n,
    a_5__n_spl_01,
    b_5__n_spl_01
  );


  and

  (
    g109_p,
    a_6__p_spl_01,
    b_3__p_spl_00
  );


  or

  (
    g109_n,
    a_6__n_spl_01,
    b_3__n_spl_00
  );


  and

  (
    g110_p,
    g17_p_spl_,
    g109_p_spl_
  );


  or

  (
    g110_n,
    g17_n_spl_,
    g109_n_spl_
  );


  and

  (
    g111_p,
    a_6__p_spl_10,
    b_4__p_spl_00
  );


  or

  (
    g111_n,
    a_6__n_spl_10,
    b_4__n_spl_00
  );


  and

  (
    g112_p,
    g19_n_spl_,
    g111_n_spl_
  );


  or

  (
    g112_n,
    g19_p_spl_,
    g111_p_spl_
  );


  and

  (
    g113_p,
    g110_n_spl_,
    g112_n
  );


  or

  (
    g113_n,
    g110_p_spl_,
    g112_p
  );


  and

  (
    g114_p,
    g108_p_spl_,
    g113_p_spl_
  );


  or

  (
    g114_n,
    g108_n_spl_,
    g113_n_spl_
  );


  and

  (
    g115_p,
    g108_n_spl_,
    g113_n_spl_
  );


  or

  (
    g115_n,
    g108_p_spl_,
    g113_p_spl_
  );


  and

  (
    g116_p,
    g114_n_spl_,
    g115_n
  );


  or

  (
    g116_n,
    g114_p_spl_,
    g115_p
  );


  and

  (
    g117_p,
    g41_p_spl_01,
    g116_p_spl_
  );


  or

  (
    g117_n,
    g41_n_spl_01,
    g116_n_spl_
  );


  and

  (
    g118_p,
    g35_n_spl_10,
    g117_n_spl_
  );


  or

  (
    g118_n,
    g35_p_spl_10,
    g117_p_spl_
  );


  and

  (
    g119_p,
    g41_n_spl_1,
    g55_n_spl_
  );


  or

  (
    g119_n,
    g41_p_spl_1,
    g55_p_spl_
  );


  and

  (
    g120_p,
    g56_n_spl_,
    g119_n
  );


  or

  (
    g120_n,
    g56_p_spl_,
    g119_p
  );


  and

  (
    g121_p,
    g118_n_spl_,
    g120_p_spl_
  );


  or

  (
    g121_n,
    g118_p_spl_,
    g120_n_spl_
  );


  and

  (
    g122_p,
    a_4__p_spl_00,
    b_6__p_spl_01
  );


  or

  (
    g122_n,
    a_4__n_spl_00,
    b_6__n_spl_01
  );


  and

  (
    g123_p,
    a_3__n_spl_00,
    b_7__p_spl_01
  );


  or

  (
    g123_n,
    a_3__p_spl_00,
    b_7__n_spl_01
  );


  and

  (
    g124_p,
    g122_p_spl_,
    g123_p_spl_
  );


  or

  (
    g124_n,
    g122_n_spl_,
    g123_n_spl_
  );


  and

  (
    g125_p,
    g110_n_spl_,
    g114_n_spl_
  );


  or

  (
    g125_n,
    g110_p_spl_,
    g114_p_spl_
  );


  and

  (
    g126_p,
    g59_n_spl_,
    g60_n_spl_
  );


  or

  (
    g126_n,
    g59_p_spl_,
    g60_p_spl_
  );


  and

  (
    g127_p,
    g61_n_spl_,
    g126_n
  );


  or

  (
    g127_n,
    g61_p_spl_,
    g126_p
  );


  and

  (
    g128_p,
    g125_n_spl_,
    g127_p_spl_
  );


  or

  (
    g128_n,
    g125_p_spl_,
    g127_n_spl_
  );


  and

  (
    g129_p,
    g125_p_spl_,
    g127_n_spl_
  );


  or

  (
    g129_n,
    g125_n_spl_,
    g127_p_spl_
  );


  and

  (
    g130_p,
    g128_n_spl_,
    g129_n
  );


  or

  (
    g130_n,
    g128_p_spl_,
    g129_p
  );


  and

  (
    g131_p,
    g124_p_spl_0,
    g130_p_spl_
  );


  or

  (
    g131_n,
    g124_n_spl_0,
    g130_n_spl_
  );


  and

  (
    g132_p,
    g124_n_spl_0,
    g130_n_spl_
  );


  or

  (
    g132_n,
    g124_p_spl_0,
    g130_p_spl_
  );


  and

  (
    g133_p,
    g131_n_spl_,
    g132_n
  );


  or

  (
    g133_n,
    g131_p_spl_,
    g132_p
  );


  and

  (
    g134_p,
    g118_p_spl_,
    g120_n_spl_
  );


  or

  (
    g134_n,
    g118_n_spl_,
    g120_p_spl_
  );


  and

  (
    g135_p,
    g121_n_spl_,
    g134_n
  );


  or

  (
    g135_n,
    g121_p_spl_,
    g134_p
  );


  and

  (
    g136_p,
    g133_p_spl_,
    g135_p_spl_
  );


  or

  (
    g136_n,
    g133_n_spl_,
    g135_n_spl_
  );


  and

  (
    g137_p,
    g121_n_spl_,
    g136_n_spl_
  );


  or

  (
    g137_n,
    g121_p_spl_,
    g136_p_spl_
  );


  and

  (
    g138_p,
    g73_n_spl_,
    g75_n_spl_
  );


  or

  (
    g138_n,
    g73_p_spl_,
    g75_p_spl_
  );


  and

  (
    g139_p,
    g76_n_spl_,
    g138_n
  );


  or

  (
    g139_n,
    g76_p_spl_,
    g138_p
  );


  and

  (
    g140_p,
    g137_n_spl_,
    g139_p_spl_
  );


  or

  (
    g140_n,
    g137_p_spl_,
    g139_n_spl_
  );


  and

  (
    g141_p,
    g128_n_spl_,
    g131_n_spl_
  );


  or

  (
    g141_n,
    g128_p_spl_,
    g131_p_spl_
  );


  and

  (
    g142_p,
    g137_p_spl_,
    g139_n_spl_
  );


  or

  (
    g142_n,
    g137_n_spl_,
    g139_p_spl_
  );


  and

  (
    g143_p,
    g140_n_spl_,
    g142_n
  );


  or

  (
    g143_n,
    g140_p_spl_,
    g142_p
  );


  and

  (
    g144_p,
    g141_n_spl_,
    g143_p_spl_
  );


  or

  (
    g144_n,
    g141_p_spl_,
    g143_n_spl_
  );


  and

  (
    g145_p,
    g140_n_spl_,
    g144_n_spl_
  );


  or

  (
    g145_n,
    g140_p_spl_,
    g144_p_spl_
  );


  and

  (
    g146_p,
    g90_p_spl_,
    g92_n_spl_
  );


  or

  (
    g146_n,
    g90_n_spl_,
    g92_p_spl_
  );


  and

  (
    g147_p,
    g93_n_spl_,
    g146_n
  );


  or

  (
    g147_n,
    g93_p_spl_,
    g146_p
  );


  and

  (
    g148_p,
    g145_n_spl_,
    g147_p_spl_
  );


  or

  (
    g148_n,
    g145_p_spl_,
    g147_n_spl_
  );


  and

  (
    g149_p,
    g145_p_spl_,
    g147_n_spl_
  );


  or

  (
    g149_n,
    g145_n_spl_,
    g147_p_spl_
  );


  and

  (
    g150_p,
    a_4__p_spl_01,
    b_5__p_spl_01
  );


  or

  (
    g150_n,
    a_4__n_spl_01,
    b_5__n_spl_01
  );


  and

  (
    g151_p,
    a_5__p_spl_01,
    b_3__p_spl_01
  );


  or

  (
    g151_n,
    a_5__n_spl_01,
    b_3__n_spl_01
  );


  and

  (
    g152_p,
    g111_p_spl_,
    g151_p_spl_0
  );


  or

  (
    g152_n,
    g111_n_spl_,
    g151_n_spl_0
  );


  and

  (
    g153_p,
    a_5__p_spl_10,
    b_4__p_spl_01
  );


  or

  (
    g153_n,
    a_5__n_spl_10,
    b_4__n_spl_01
  );


  and

  (
    g154_p,
    g109_n_spl_,
    g153_n
  );


  or

  (
    g154_n,
    g109_p_spl_,
    g153_p
  );


  and

  (
    g155_p,
    g152_n_spl_,
    g154_n
  );


  or

  (
    g155_n,
    g152_p_spl_,
    g154_p
  );


  and

  (
    g156_p,
    g150_p_spl_,
    g155_p_spl_
  );


  or

  (
    g156_n,
    g150_n_spl_,
    g155_n_spl_
  );


  and

  (
    g157_p,
    g150_n_spl_,
    g155_n_spl_
  );


  or

  (
    g157_n,
    g150_p_spl_,
    g155_p_spl_
  );


  and

  (
    g158_p,
    g156_n_spl_,
    g157_n
  );


  or

  (
    g158_n,
    g156_p_spl_,
    g157_p
  );


  and

  (
    g159_p,
    a_6__p_spl_10,
    b_2__p_spl_00
  );


  or

  (
    g159_n,
    a_6__n_spl_10,
    b_2__n_spl_00
  );


  and

  (
    g160_p,
    g37_p_spl_,
    g159_n_spl_0
  );


  or

  (
    g160_n,
    g37_n_spl_,
    g159_p_spl_0
  );


  and

  (
    g161_p,
    g39_p_spl_0,
    g160_p
  );


  or

  (
    g161_n,
    g39_n_spl_0,
    g160_n
  );


  and

  (
    g162_p,
    g40_n_spl_,
    g161_n
  );


  or

  (
    g162_n,
    g40_p_spl_,
    g161_p
  );


  and

  (
    g163_p,
    g34_n_spl_0,
    g162_n
  );


  or

  (
    g163_n,
    g34_p_spl_0,
    g162_p
  );


  and

  (
    g164_p,
    g35_n_spl_10,
    g163_n
  );


  or

  (
    g164_n,
    g35_p_spl_10,
    g163_p
  );


  and

  (
    g165_p,
    g158_p_spl_,
    g164_p_spl_
  );


  or

  (
    g165_n,
    g158_n_spl_,
    g164_n_spl_
  );


  and

  (
    g166_p,
    g35_n_spl_1,
    g165_n_spl_
  );


  or

  (
    g166_n,
    g35_p_spl_1,
    g165_p_spl_
  );


  and

  (
    g167_p,
    g41_n_spl_1,
    g116_n_spl_
  );


  or

  (
    g167_n,
    g41_p_spl_1,
    g116_p_spl_
  );


  and

  (
    g168_p,
    g117_n_spl_,
    g167_n
  );


  or

  (
    g168_n,
    g117_p_spl_,
    g167_p
  );


  and

  (
    g169_p,
    g166_n_spl_,
    g168_p_spl_
  );


  or

  (
    g169_n,
    g166_p_spl_,
    g168_n_spl_
  );


  and

  (
    g170_p,
    a_3__p_spl_00,
    b_6__p_spl_10
  );


  or

  (
    g170_n,
    a_3__n_spl_00,
    b_6__n_spl_10
  );


  and

  (
    g171_p,
    a_2__n_spl_00,
    b_7__p_spl_01
  );


  or

  (
    g171_n,
    a_2__p_spl_00,
    b_7__n_spl_01
  );


  and

  (
    g172_p,
    g170_p_spl_,
    g171_p_spl_
  );


  or

  (
    g172_n,
    g170_n_spl_,
    g171_n_spl_
  );


  and

  (
    g173_p,
    g152_n_spl_,
    g156_n_spl_
  );


  or

  (
    g173_n,
    g152_p_spl_,
    g156_p_spl_
  );


  and

  (
    g174_p,
    g122_n_spl_,
    g123_n_spl_
  );


  or

  (
    g174_n,
    g122_p_spl_,
    g123_p_spl_
  );


  and

  (
    g175_p,
    g124_n_spl_,
    g174_n
  );


  or

  (
    g175_n,
    g124_p_spl_,
    g174_p
  );


  and

  (
    g176_p,
    g173_n_spl_,
    g175_p_spl_
  );


  or

  (
    g176_n,
    g173_p_spl_,
    g175_n_spl_
  );


  and

  (
    g177_p,
    g173_p_spl_,
    g175_n_spl_
  );


  or

  (
    g177_n,
    g173_n_spl_,
    g175_p_spl_
  );


  and

  (
    g178_p,
    g176_n_spl_,
    g177_n
  );


  or

  (
    g178_n,
    g176_p_spl_,
    g177_p
  );


  and

  (
    g179_p,
    g172_p_spl_0,
    g178_p_spl_
  );


  or

  (
    g179_n,
    g172_n_spl_0,
    g178_n_spl_
  );


  and

  (
    g180_p,
    g172_n_spl_0,
    g178_n_spl_
  );


  or

  (
    g180_n,
    g172_p_spl_0,
    g178_p_spl_
  );


  and

  (
    g181_p,
    g179_n_spl_,
    g180_n
  );


  or

  (
    g181_n,
    g179_p_spl_,
    g180_p
  );


  and

  (
    g182_p,
    g166_p_spl_,
    g168_n_spl_
  );


  or

  (
    g182_n,
    g166_n_spl_,
    g168_p_spl_
  );


  and

  (
    g183_p,
    g169_n_spl_,
    g182_n
  );


  or

  (
    g183_n,
    g169_p_spl_,
    g182_p
  );


  and

  (
    g184_p,
    g181_p_spl_,
    g183_p_spl_
  );


  or

  (
    g184_n,
    g181_n_spl_,
    g183_n_spl_
  );


  and

  (
    g185_p,
    g169_n_spl_,
    g184_n_spl_
  );


  or

  (
    g185_n,
    g169_p_spl_,
    g184_p_spl_
  );


  and

  (
    g186_p,
    g133_n_spl_,
    g135_n_spl_
  );


  or

  (
    g186_n,
    g133_p_spl_,
    g135_p_spl_
  );


  and

  (
    g187_p,
    g136_n_spl_,
    g186_n
  );


  or

  (
    g187_n,
    g136_p_spl_,
    g186_p
  );


  and

  (
    g188_p,
    g185_n_spl_,
    g187_p_spl_
  );


  or

  (
    g188_n,
    g185_p_spl_,
    g187_n_spl_
  );


  and

  (
    g189_p,
    g176_n_spl_,
    g179_n_spl_
  );


  or

  (
    g189_n,
    g176_p_spl_,
    g179_p_spl_
  );


  and

  (
    g190_p,
    g185_p_spl_,
    g187_n_spl_
  );


  or

  (
    g190_n,
    g185_n_spl_,
    g187_p_spl_
  );


  and

  (
    g191_p,
    g188_n_spl_,
    g190_n
  );


  or

  (
    g191_n,
    g188_p_spl_,
    g190_p
  );


  and

  (
    g192_p,
    g189_n_spl_,
    g191_p_spl_
  );


  or

  (
    g192_n,
    g189_p_spl_,
    g191_n_spl_
  );


  and

  (
    g193_p,
    g188_n_spl_,
    g192_n_spl_
  );


  or

  (
    g193_n,
    g188_p_spl_,
    g192_p_spl_
  );


  and

  (
    g194_p,
    g141_p_spl_,
    g143_n_spl_
  );


  or

  (
    g194_n,
    g141_n_spl_,
    g143_p_spl_
  );


  and

  (
    g195_p,
    g144_n_spl_,
    g194_n
  );


  or

  (
    g195_n,
    g144_p_spl_,
    g194_p
  );


  and

  (
    g196_p,
    g193_n_spl_,
    g195_p_spl_
  );


  or

  (
    g196_n,
    g193_p_spl_,
    g195_n_spl_
  );


  and

  (
    g197_p,
    b_7__p_spl_10,
    g33_p_spl_0
  );


  or

  (
    g197_n,
    b_7__n_spl_10,
    g33_n_spl_0
  );


  and

  (
    g198_p,
    a_6__p_spl_11,
    b_1__p_spl_00
  );


  or

  (
    g198_n,
    a_6__n_spl_11,
    b_1__n_spl_01
  );


  and

  (
    g199_p,
    b_7__n_spl_10,
    g33_n_spl_
  );


  or

  (
    g199_n,
    b_7__p_spl_10,
    g33_p_spl_
  );


  and

  (
    g200_p,
    g197_n_spl_,
    g199_n
  );


  or

  (
    g200_n,
    g197_p_spl_,
    g199_p
  );


  and

  (
    g201_p,
    g198_p_spl_0,
    g200_p_spl_
  );


  or

  (
    g201_n,
    g198_n_spl_0,
    g200_n_spl_
  );


  and

  (
    g202_p,
    g197_n_spl_,
    g201_n_spl_
  );


  or

  (
    g202_n,
    g197_p_spl_,
    g201_p_spl_
  );


  and

  (
    g203_p,
    g34_n_spl_,
    g39_p_spl_
  );


  or

  (
    g203_n,
    g34_p_spl_,
    g39_n_spl_
  );


  and

  (
    g204_p,
    g159_n_spl_0,
    g203_p_spl_
  );


  or

  (
    g204_n,
    g159_p_spl_0,
    g203_n_spl_
  );


  and

  (
    g205_p,
    g159_p_spl_,
    g203_n_spl_
  );


  or

  (
    g205_n,
    g159_n_spl_,
    g203_p_spl_
  );


  and

  (
    g206_p,
    g204_n,
    g205_n
  );


  or

  (
    g206_n,
    g204_p,
    g205_p
  );


  and

  (
    g207_p,
    g202_n_spl_,
    g206_n_spl_
  );


  or

  (
    g207_n,
    g202_p_spl_,
    g206_p_spl_
  );


  and

  (
    g208_p,
    a_3__p_spl_01,
    b_5__p_spl_10
  );


  or

  (
    g208_n,
    a_3__n_spl_01,
    b_5__n_spl_10
  );


  and

  (
    g209_p,
    a_4__p_spl_01,
    b_4__p_spl_01
  );


  or

  (
    g209_n,
    a_4__n_spl_01,
    b_4__n_spl_01
  );


  and

  (
    g210_p,
    g151_p_spl_0,
    g209_p_spl_
  );


  or

  (
    g210_n,
    g151_n_spl_0,
    g209_n_spl_
  );


  and

  (
    g211_p,
    g151_n_spl_1,
    g209_n_spl_
  );


  or

  (
    g211_n,
    g151_p_spl_1,
    g209_p_spl_
  );


  and

  (
    g212_p,
    g210_n_spl_,
    g211_n
  );


  or

  (
    g212_n,
    g210_p_spl_,
    g211_p
  );


  and

  (
    g213_p,
    g208_p_spl_,
    g212_p_spl_
  );


  or

  (
    g213_n,
    g208_n_spl_,
    g212_n_spl_
  );


  and

  (
    g214_p,
    g208_n_spl_,
    g212_n_spl_
  );


  or

  (
    g214_n,
    g208_p_spl_,
    g212_p_spl_
  );


  and

  (
    g215_p,
    g213_n_spl_,
    g214_n
  );


  or

  (
    g215_n,
    g213_p_spl_,
    g214_p
  );


  and

  (
    g216_p,
    g202_p_spl_,
    g206_p_spl_
  );


  or

  (
    g216_n,
    g202_n_spl_,
    g206_n_spl_
  );


  and

  (
    g217_p,
    g207_n_spl_,
    g216_n
  );


  or

  (
    g217_n,
    g207_p_spl_,
    g216_p
  );


  and

  (
    g218_p,
    g215_p_spl_,
    g217_p_spl_
  );


  or

  (
    g218_n,
    g215_n_spl_,
    g217_n_spl_
  );


  and

  (
    g219_p,
    g207_n_spl_,
    g218_n_spl_
  );


  or

  (
    g219_n,
    g207_p_spl_,
    g218_p_spl_
  );


  and

  (
    g220_p,
    g158_n_spl_,
    g164_n_spl_
  );


  or

  (
    g220_n,
    g158_p_spl_,
    g164_p_spl_
  );


  and

  (
    g221_p,
    g165_n_spl_,
    g220_n
  );


  or

  (
    g221_n,
    g165_p_spl_,
    g220_p
  );


  and

  (
    g222_p,
    g219_n_spl_,
    g221_p_spl_
  );


  or

  (
    g222_n,
    g219_p_spl_,
    g221_n_spl_
  );


  and

  (
    g223_p,
    a_2__p_spl_00,
    b_6__p_spl_10
  );


  or

  (
    g223_n,
    a_2__n_spl_00,
    b_6__n_spl_10
  );


  and

  (
    g224_p,
    a_1__n_spl_00,
    b_7__p_spl_11
  );


  or

  (
    g224_n,
    a_1__p_spl_00,
    b_7__n_spl_11
  );


  and

  (
    g225_p,
    g223_p_spl_0,
    g224_p_spl_
  );


  or

  (
    g225_n,
    g223_n_spl_0,
    g224_n_spl_
  );


  and

  (
    g226_p,
    g210_n_spl_,
    g213_n_spl_
  );


  or

  (
    g226_n,
    g210_p_spl_,
    g213_p_spl_
  );


  and

  (
    g227_p,
    g170_n_spl_,
    g171_n_spl_
  );


  or

  (
    g227_n,
    g170_p_spl_,
    g171_p_spl_
  );


  and

  (
    g228_p,
    g172_n_spl_,
    g227_n
  );


  or

  (
    g228_n,
    g172_p_spl_,
    g227_p
  );


  and

  (
    g229_p,
    g226_n_spl_,
    g228_p_spl_
  );


  or

  (
    g229_n,
    g226_p_spl_,
    g228_n_spl_
  );


  and

  (
    g230_p,
    g226_p_spl_,
    g228_n_spl_
  );


  or

  (
    g230_n,
    g226_n_spl_,
    g228_p_spl_
  );


  and

  (
    g231_p,
    g229_n_spl_,
    g230_n
  );


  or

  (
    g231_n,
    g229_p_spl_,
    g230_p
  );


  and

  (
    g232_p,
    g225_p_spl_0,
    g231_p_spl_
  );


  or

  (
    g232_n,
    g225_n_spl_0,
    g231_n_spl_
  );


  and

  (
    g233_p,
    g225_n_spl_0,
    g231_n_spl_
  );


  or

  (
    g233_n,
    g225_p_spl_0,
    g231_p_spl_
  );


  and

  (
    g234_p,
    g232_n_spl_,
    g233_n
  );


  or

  (
    g234_n,
    g232_p_spl_,
    g233_p
  );


  and

  (
    g235_p,
    g219_p_spl_,
    g221_n_spl_
  );


  or

  (
    g235_n,
    g219_n_spl_,
    g221_p_spl_
  );


  and

  (
    g236_p,
    g222_n_spl_,
    g235_n
  );


  or

  (
    g236_n,
    g222_p_spl_,
    g235_p
  );


  and

  (
    g237_p,
    g234_p_spl_,
    g236_p_spl_
  );


  or

  (
    g237_n,
    g234_n_spl_,
    g236_n_spl_
  );


  and

  (
    g238_p,
    g222_n_spl_,
    g237_n_spl_
  );


  or

  (
    g238_n,
    g222_p_spl_,
    g237_p_spl_
  );


  and

  (
    g239_p,
    g181_n_spl_,
    g183_n_spl_
  );


  or

  (
    g239_n,
    g181_p_spl_,
    g183_p_spl_
  );


  and

  (
    g240_p,
    g184_n_spl_,
    g239_n
  );


  or

  (
    g240_n,
    g184_p_spl_,
    g239_p
  );


  and

  (
    g241_p,
    g238_n_spl_,
    g240_p_spl_
  );


  or

  (
    g241_n,
    g238_p_spl_,
    g240_n_spl_
  );


  and

  (
    g242_p,
    g229_n_spl_,
    g232_n_spl_
  );


  or

  (
    g242_n,
    g229_p_spl_,
    g232_p_spl_
  );


  and

  (
    g243_p,
    g238_p_spl_,
    g240_n_spl_
  );


  or

  (
    g243_n,
    g238_n_spl_,
    g240_p_spl_
  );


  and

  (
    g244_p,
    g241_n_spl_,
    g243_n
  );


  or

  (
    g244_n,
    g241_p_spl_,
    g243_p
  );


  and

  (
    g245_p,
    g242_n_spl_,
    g244_p_spl_
  );


  or

  (
    g245_n,
    g242_p_spl_,
    g244_n_spl_
  );


  and

  (
    g246_p,
    g241_n_spl_,
    g245_n_spl_
  );


  or

  (
    g246_n,
    g241_p_spl_,
    g245_p_spl_
  );


  and

  (
    g247_p,
    g189_p_spl_,
    g191_n_spl_
  );


  or

  (
    g247_n,
    g189_n_spl_,
    g191_p_spl_
  );


  and

  (
    g248_p,
    g192_n_spl_,
    g247_n
  );


  or

  (
    g248_n,
    g192_p_spl_,
    g247_p
  );


  and

  (
    g249_p,
    g246_n_spl_,
    g248_p_spl_
  );


  or

  (
    g249_n,
    g246_p_spl_,
    g248_n_spl_
  );


  and

  (
    g250_p,
    g246_p_spl_,
    g248_n_spl_
  );


  or

  (
    g250_n,
    g246_n_spl_,
    g248_p_spl_
  );


  and

  (
    g251_p,
    g249_n_spl_,
    g250_n
  );


  or

  (
    g251_n,
    g249_p_spl_,
    g250_p
  );


  and

  (
    g252_p,
    a_5__p_spl_10,
    b_0__p_spl_00
  );


  or

  (
    g252_n,
    a_5__n_spl_10,
    b_0__n_spl_01
  );


  and

  (
    g253_p,
    g198_p_spl_0,
    g252_p_spl_0
  );


  or

  (
    g253_n,
    g198_n_spl_0,
    g252_n_spl_0
  );


  and

  (
    g254_p,
    a_4__p_spl_10,
    b_2__p_spl_01
  );


  or

  (
    g254_n,
    a_4__n_spl_10,
    b_2__n_spl_01
  );


  and

  (
    g255_p,
    a_6__p_spl_11,
    b_0__p_spl_01
  );


  or

  (
    g255_n,
    a_6__n_spl_11,
    b_0__n_spl_01
  );


  and

  (
    g256_p,
    a_5__p_spl_11,
    b_1__p_spl_01
  );


  or

  (
    g256_n,
    a_5__n_spl_11,
    b_1__n_spl_01
  );


  and

  (
    g257_p,
    g255_n,
    g256_n
  );


  or

  (
    g257_n,
    g255_p,
    g256_p
  );


  and

  (
    g258_p,
    g253_n_spl_,
    g257_n
  );


  or

  (
    g258_n,
    g253_p_spl_,
    g257_p
  );


  and

  (
    g259_p,
    g254_p_spl_0,
    g258_p_spl_
  );


  or

  (
    g259_n,
    g254_n_spl_0,
    g258_n_spl_
  );


  and

  (
    g260_p,
    g253_n_spl_,
    g259_n_spl_
  );


  or

  (
    g260_n,
    g253_p_spl_,
    g259_p_spl_
  );


  and

  (
    g261_p,
    g198_n_spl_,
    g200_n_spl_
  );


  or

  (
    g261_n,
    g198_p_spl_,
    g200_p_spl_
  );


  and

  (
    g262_p,
    g201_n_spl_,
    g261_n
  );


  or

  (
    g262_n,
    g201_p_spl_,
    g261_p
  );


  and

  (
    g263_p,
    g260_n_spl_,
    g262_p_spl_
  );


  or

  (
    g263_n,
    g260_p_spl_,
    g262_n_spl_
  );


  and

  (
    g264_p,
    a_3__p_spl_01,
    b_4__p_spl_10
  );


  or

  (
    g264_n,
    a_3__n_spl_01,
    b_4__n_spl_10
  );


  and

  (
    g265_p,
    g151_p_spl_1,
    g254_p_spl_0
  );


  or

  (
    g265_n,
    g151_n_spl_1,
    g254_n_spl_0
  );


  and

  (
    g266_p,
    a_4__p_spl_10,
    b_3__p_spl_01
  );


  or

  (
    g266_n,
    a_4__n_spl_10,
    b_3__n_spl_01
  );


  and

  (
    g267_p,
    a_5__p_spl_11,
    b_2__p_spl_01
  );


  or

  (
    g267_n,
    a_5__n_spl_11,
    b_2__n_spl_01
  );


  and

  (
    g268_p,
    g266_n,
    g267_n
  );


  or

  (
    g268_n,
    g266_p,
    g267_p
  );


  and

  (
    g269_p,
    g265_n_spl_,
    g268_n
  );


  or

  (
    g269_n,
    g265_p_spl_,
    g268_p
  );


  and

  (
    g270_p,
    g264_p_spl_0,
    g269_p_spl_
  );


  or

  (
    g270_n,
    g264_n_spl_0,
    g269_n_spl_
  );


  and

  (
    g271_p,
    g264_n_spl_0,
    g269_n_spl_
  );


  or

  (
    g271_n,
    g264_p_spl_0,
    g269_p_spl_
  );


  and

  (
    g272_p,
    g270_n_spl_,
    g271_n
  );


  or

  (
    g272_n,
    g270_p_spl_,
    g271_p
  );


  and

  (
    g273_p,
    g260_p_spl_,
    g262_n_spl_
  );


  or

  (
    g273_n,
    g260_n_spl_,
    g262_p_spl_
  );


  and

  (
    g274_p,
    g263_n_spl_,
    g273_n
  );


  or

  (
    g274_n,
    g263_p_spl_,
    g273_p
  );


  and

  (
    g275_p,
    g272_p_spl_,
    g274_p_spl_
  );


  or

  (
    g275_n,
    g272_n_spl_,
    g274_n_spl_
  );


  and

  (
    g276_p,
    g263_n_spl_,
    g275_n_spl_
  );


  or

  (
    g276_n,
    g263_p_spl_,
    g275_p_spl_
  );


  and

  (
    g277_p,
    g215_n_spl_,
    g217_n_spl_
  );


  or

  (
    g277_n,
    g215_p_spl_,
    g217_p_spl_
  );


  and

  (
    g278_p,
    g218_n_spl_,
    g277_n
  );


  or

  (
    g278_n,
    g218_p_spl_,
    g277_p
  );


  and

  (
    g279_p,
    g276_n_spl_,
    g278_p_spl_
  );


  or

  (
    g279_n,
    g276_p_spl_,
    g278_n_spl_
  );


  and

  (
    g280_p,
    a_1__p_spl_00,
    b_5__p_spl_10
  );


  or

  (
    g280_n,
    a_1__n_spl_00,
    b_5__n_spl_10
  );


  and

  (
    g281_p,
    g223_p_spl_0,
    g280_p_spl_0
  );


  or

  (
    g281_n,
    g223_n_spl_0,
    g280_n_spl_0
  );


  and

  (
    g282_p,
    a_0__n_spl_00,
    b_7__p_spl_11
  );


  or

  (
    g282_n,
    a_0__p_spl_00,
    b_7__n_spl_11
  );


  and

  (
    g283_p,
    a_2__p_spl_01,
    b_5__p_spl_11
  );


  or

  (
    g283_n,
    a_2__n_spl_01,
    b_5__n_spl_11
  );


  and

  (
    g284_p,
    a_1__p_spl_01,
    b_6__p_spl_11
  );


  or

  (
    g284_n,
    a_1__n_spl_01,
    b_6__n_spl_11
  );


  and

  (
    g285_p,
    g283_n,
    g284_n
  );


  or

  (
    g285_n,
    g283_p,
    g284_p
  );


  and

  (
    g286_p,
    g281_n_spl_,
    g285_n
  );


  or

  (
    g286_n,
    g281_p_spl_,
    g285_p
  );


  and

  (
    g287_p,
    g282_p_spl_,
    g286_p_spl_
  );


  or

  (
    g287_n,
    g282_n_spl_,
    g286_n_spl_
  );


  and

  (
    g288_p,
    g281_n_spl_,
    g287_n_spl_
  );


  or

  (
    g288_n,
    g281_p_spl_,
    g287_p_spl_
  );


  and

  (
    g289_p,
    g265_n_spl_,
    g270_n_spl_
  );


  or

  (
    g289_n,
    g265_p_spl_,
    g270_p_spl_
  );


  and

  (
    g290_p,
    g223_n_spl_,
    g224_n_spl_
  );


  or

  (
    g290_n,
    g223_p_spl_,
    g224_p_spl_
  );


  and

  (
    g291_p,
    g225_n_spl_,
    g290_n
  );


  or

  (
    g291_n,
    g225_p_spl_,
    g290_p
  );


  and

  (
    g292_p,
    g289_n_spl_,
    g291_p_spl_
  );


  or

  (
    g292_n,
    g289_p_spl_,
    g291_n_spl_
  );


  and

  (
    g293_p,
    g289_p_spl_,
    g291_n_spl_
  );


  or

  (
    g293_n,
    g289_n_spl_,
    g291_p_spl_
  );


  and

  (
    g294_p,
    g292_n_spl_,
    g293_n
  );


  or

  (
    g294_n,
    g292_p_spl_,
    g293_p
  );


  and

  (
    g295_p,
    g288_n_spl_,
    g294_p_spl_
  );


  or

  (
    g295_n,
    g288_p_spl_,
    g294_n_spl_
  );


  and

  (
    g296_p,
    g288_p_spl_,
    g294_n_spl_
  );


  or

  (
    g296_n,
    g288_n_spl_,
    g294_p_spl_
  );


  and

  (
    g297_p,
    g295_n_spl_,
    g296_n
  );


  or

  (
    g297_n,
    g295_p_spl_,
    g296_p
  );


  and

  (
    g298_p,
    g276_p_spl_,
    g278_n_spl_
  );


  or

  (
    g298_n,
    g276_n_spl_,
    g278_p_spl_
  );


  and

  (
    g299_p,
    g279_n_spl_,
    g298_n
  );


  or

  (
    g299_n,
    g279_p_spl_,
    g298_p
  );


  and

  (
    g300_p,
    g297_p_spl_,
    g299_p_spl_
  );


  or

  (
    g300_n,
    g297_n_spl_,
    g299_n_spl_
  );


  and

  (
    g301_p,
    g279_n_spl_,
    g300_n_spl_
  );


  or

  (
    g301_n,
    g279_p_spl_,
    g300_p_spl_
  );


  and

  (
    g302_p,
    g234_n_spl_,
    g236_n_spl_
  );


  or

  (
    g302_n,
    g234_p_spl_,
    g236_p_spl_
  );


  and

  (
    g303_p,
    g237_n_spl_,
    g302_n
  );


  or

  (
    g303_n,
    g237_p_spl_,
    g302_p
  );


  and

  (
    g304_p,
    g301_n_spl_,
    g303_p_spl_
  );


  or

  (
    g304_n,
    g301_p_spl_,
    g303_n_spl_
  );


  and

  (
    g305_p,
    g292_n_spl_,
    g295_n_spl_
  );


  or

  (
    g305_n,
    g292_p_spl_,
    g295_p_spl_
  );


  and

  (
    g306_p,
    g301_p_spl_,
    g303_n_spl_
  );


  or

  (
    g306_n,
    g301_n_spl_,
    g303_p_spl_
  );


  and

  (
    g307_p,
    g304_n_spl_,
    g306_n
  );


  or

  (
    g307_n,
    g304_p_spl_,
    g306_p
  );


  and

  (
    g308_p,
    g305_n_spl_,
    g307_p_spl_
  );


  or

  (
    g308_n,
    g305_p_spl_,
    g307_n_spl_
  );


  and

  (
    g309_p,
    g304_n_spl_,
    g308_n_spl_
  );


  or

  (
    g309_n,
    g304_p_spl_,
    g308_p_spl_
  );


  and

  (
    g310_p,
    g242_p_spl_,
    g244_n_spl_
  );


  or

  (
    g310_n,
    g242_n_spl_,
    g244_p_spl_
  );


  and

  (
    g311_p,
    g245_n_spl_,
    g310_n
  );


  or

  (
    g311_n,
    g245_p_spl_,
    g310_p
  );


  and

  (
    g312_p,
    g309_n_spl_,
    g311_p_spl_
  );


  or

  (
    g312_n,
    g309_p_spl_,
    g311_n_spl_
  );


  and

  (
    g313_p,
    g309_p_spl_,
    g311_n_spl_
  );


  or

  (
    g313_n,
    g309_n_spl_,
    g311_p_spl_
  );


  and

  (
    g314_p,
    g312_n_spl_,
    g313_n
  );


  or

  (
    g314_n,
    g312_p_spl_,
    g313_p
  );


  and

  (
    g315_p,
    a_4__p_spl_11,
    b_1__p_spl_01
  );


  or

  (
    g315_n,
    a_4__n_spl_11,
    b_1__n_spl_10
  );


  and

  (
    g316_p,
    g252_p_spl_0,
    g315_p_spl_
  );


  or

  (
    g316_n,
    g252_n_spl_0,
    g315_n_spl_
  );


  and

  (
    g317_p,
    a_3__p_spl_10,
    b_2__p_spl_10
  );


  or

  (
    g317_n,
    a_3__n_spl_10,
    b_2__n_spl_10
  );


  and

  (
    g318_p,
    g252_n_spl_,
    g315_n_spl_
  );


  or

  (
    g318_n,
    g252_p_spl_,
    g315_p_spl_
  );


  and

  (
    g319_p,
    g316_n_spl_,
    g318_n
  );


  or

  (
    g319_n,
    g316_p_spl_,
    g318_p
  );


  and

  (
    g320_p,
    g317_p_spl_,
    g319_p_spl_
  );


  or

  (
    g320_n,
    g317_n_spl_,
    g319_n_spl_
  );


  and

  (
    g321_p,
    g316_n_spl_,
    g320_n_spl_
  );


  or

  (
    g321_n,
    g316_p_spl_,
    g320_p_spl_
  );


  and

  (
    g322_p,
    g254_n_spl_,
    g258_n_spl_
  );


  or

  (
    g322_n,
    g254_p_spl_,
    g258_p_spl_
  );


  and

  (
    g323_p,
    g259_n_spl_,
    g322_n
  );


  or

  (
    g323_n,
    g259_p_spl_,
    g322_p
  );


  and

  (
    g324_p,
    g321_n_spl_,
    g323_p_spl_
  );


  or

  (
    g324_n,
    g321_p_spl_,
    g323_n_spl_
  );


  and

  (
    g325_p,
    a_2__p_spl_01,
    b_3__p_spl_10
  );


  or

  (
    g325_n,
    a_2__n_spl_01,
    b_3__n_spl_10
  );


  and

  (
    g326_p,
    g264_p_spl_,
    g325_p_spl_0
  );


  or

  (
    g326_n,
    g264_n_spl_,
    g325_n_spl_0
  );


  and

  (
    g327_p,
    a_3__p_spl_10,
    b_3__p_spl_10
  );


  or

  (
    g327_n,
    a_3__n_spl_10,
    b_3__n_spl_10
  );


  and

  (
    g328_p,
    a_2__p_spl_10,
    b_4__p_spl_10
  );


  or

  (
    g328_n,
    a_2__n_spl_10,
    b_4__n_spl_10
  );


  and

  (
    g329_p,
    g327_n,
    g328_n
  );


  or

  (
    g329_n,
    g327_p,
    g328_p
  );


  and

  (
    g330_p,
    g326_n_spl_,
    g329_n
  );


  or

  (
    g330_n,
    g326_p_spl_,
    g329_p
  );


  and

  (
    g331_p,
    g280_p_spl_0,
    g330_p_spl_
  );


  or

  (
    g331_n,
    g280_n_spl_0,
    g330_n_spl_
  );


  and

  (
    g332_p,
    g280_n_spl_,
    g330_n_spl_
  );


  or

  (
    g332_n,
    g280_p_spl_,
    g330_p_spl_
  );


  and

  (
    g333_p,
    g331_n_spl_,
    g332_n
  );


  or

  (
    g333_n,
    g331_p_spl_,
    g332_p
  );


  and

  (
    g334_p,
    g321_p_spl_,
    g323_n_spl_
  );


  or

  (
    g334_n,
    g321_n_spl_,
    g323_p_spl_
  );


  and

  (
    g335_p,
    g324_n_spl_,
    g334_n
  );


  or

  (
    g335_n,
    g324_p_spl_,
    g334_p
  );


  and

  (
    g336_p,
    g333_p_spl_,
    g335_p_spl_
  );


  or

  (
    g336_n,
    g333_n_spl_,
    g335_n_spl_
  );


  and

  (
    g337_p,
    g324_n_spl_,
    g336_n_spl_
  );


  or

  (
    g337_n,
    g324_p_spl_,
    g336_p_spl_
  );


  and

  (
    g338_p,
    g272_n_spl_,
    g274_n_spl_
  );


  or

  (
    g338_n,
    g272_p_spl_,
    g274_p_spl_
  );


  and

  (
    g339_p,
    g275_n_spl_,
    g338_n
  );


  or

  (
    g339_n,
    g275_p_spl_,
    g338_p
  );


  and

  (
    g340_p,
    g337_n_spl_,
    g339_p_spl_
  );


  or

  (
    g340_n,
    g337_p_spl_,
    g339_n_spl_
  );


  and

  (
    g341_p,
    g326_n_spl_,
    g331_n_spl_
  );


  or

  (
    g341_n,
    g326_p_spl_,
    g331_p_spl_
  );


  and

  (
    g342_p,
    g282_n_spl_,
    g286_n_spl_
  );


  or

  (
    g342_n,
    g282_p_spl_,
    g286_p_spl_
  );


  and

  (
    g343_p,
    g287_n_spl_,
    g342_n
  );


  or

  (
    g343_n,
    g287_p_spl_,
    g342_p
  );


  and

  (
    g344_p,
    g341_n_spl_,
    g343_p_spl_
  );


  or

  (
    g344_n,
    g341_p_spl_,
    g343_n_spl_
  );


  and

  (
    g345_p,
    g341_p_spl_,
    g343_n_spl_
  );


  or

  (
    g345_n,
    g341_n_spl_,
    g343_p_spl_
  );


  and

  (
    g346_p,
    g344_n_spl_0,
    g345_n
  );


  or

  (
    g346_n,
    g344_p_spl_0,
    g345_p
  );


  and

  (
    g347_p,
    g337_p_spl_,
    g339_n_spl_
  );


  or

  (
    g347_n,
    g337_n_spl_,
    g339_p_spl_
  );


  and

  (
    g348_p,
    g340_n_spl_,
    g347_n
  );


  or

  (
    g348_n,
    g340_p_spl_,
    g347_p
  );


  and

  (
    g349_p,
    g346_p_spl_,
    g348_p_spl_
  );


  or

  (
    g349_n,
    g346_n_spl_,
    g348_n_spl_
  );


  and

  (
    g350_p,
    g340_n_spl_,
    g349_n_spl_
  );


  or

  (
    g350_n,
    g340_p_spl_,
    g349_p_spl_
  );


  and

  (
    g351_p,
    g297_n_spl_,
    g299_n_spl_
  );


  or

  (
    g351_n,
    g297_p_spl_,
    g299_p_spl_
  );


  and

  (
    g352_p,
    g300_n_spl_,
    g351_n
  );


  or

  (
    g352_n,
    g300_p_spl_,
    g351_p
  );


  and

  (
    g353_p,
    g350_n_spl_,
    g352_p_spl_
  );


  or

  (
    g353_n,
    g350_p_spl_,
    g352_n_spl_
  );


  and

  (
    g354_p,
    g350_p_spl_,
    g352_n_spl_
  );


  or

  (
    g354_n,
    g350_n_spl_,
    g352_p_spl_
  );


  and

  (
    g355_p,
    g353_n_spl_,
    g354_n
  );


  or

  (
    g355_n,
    g353_p_spl_,
    g354_p
  );


  and

  (
    g356_p,
    g344_p_spl_0,
    g355_p_spl_
  );


  or

  (
    g356_n,
    g344_n_spl_0,
    g355_n_spl_
  );


  and

  (
    g357_p,
    g353_n_spl_,
    g356_n_spl_
  );


  or

  (
    g357_n,
    g353_p_spl_,
    g356_p_spl_
  );


  and

  (
    g358_p,
    g305_p_spl_,
    g307_n_spl_
  );


  or

  (
    g358_n,
    g305_n_spl_,
    g307_p_spl_
  );


  and

  (
    g359_p,
    g308_n_spl_,
    g358_n
  );


  or

  (
    g359_n,
    g308_p_spl_,
    g358_p
  );


  and

  (
    g360_p,
    g357_n_spl_,
    g359_p_spl_
  );


  or

  (
    g360_n,
    g357_p_spl_,
    g359_n_spl_
  );


  and

  (
    g361_p,
    a_4__p_spl_11,
    b_0__p_spl_01
  );


  or

  (
    g361_n,
    a_4__n_spl_11,
    b_0__n_spl_10
  );


  and

  (
    g362_p,
    a_3__p_spl_11,
    b_1__p_spl_10
  );


  or

  (
    g362_n,
    a_3__n_spl_11,
    b_1__n_spl_10
  );


  and

  (
    g363_p,
    g361_p_spl_,
    g362_p_spl_0
  );


  or

  (
    g363_n,
    g361_n_spl_,
    g362_n_spl_0
  );


  and

  (
    g364_p,
    a_2__p_spl_10,
    b_2__p_spl_10
  );


  or

  (
    g364_n,
    a_2__n_spl_10,
    b_2__n_spl_10
  );


  and

  (
    g365_p,
    g361_n_spl_,
    g362_n_spl_0
  );


  or

  (
    g365_n,
    g361_p_spl_,
    g362_p_spl_0
  );


  and

  (
    g366_p,
    g363_n_spl_,
    g365_n
  );


  or

  (
    g366_n,
    g363_p_spl_,
    g365_p
  );


  and

  (
    g367_p,
    g364_p_spl_,
    g366_p_spl_
  );


  or

  (
    g367_n,
    g364_n_spl_,
    g366_n_spl_
  );


  and

  (
    g368_p,
    g363_n_spl_,
    g367_n_spl_
  );


  or

  (
    g368_n,
    g363_p_spl_,
    g367_p_spl_
  );


  and

  (
    g369_p,
    g317_n_spl_,
    g319_n_spl_
  );


  or

  (
    g369_n,
    g317_p_spl_,
    g319_p_spl_
  );


  and

  (
    g370_p,
    g320_n_spl_,
    g369_n
  );


  or

  (
    g370_n,
    g320_p_spl_,
    g369_p
  );


  and

  (
    g371_p,
    g368_n_spl_,
    g370_p_spl_
  );


  or

  (
    g371_n,
    g368_p_spl_,
    g370_n_spl_
  );


  and

  (
    g372_p,
    a_0__p_spl_00,
    b_5__p_spl_11
  );


  or

  (
    g372_n,
    a_0__n_spl_00,
    b_5__n_spl_11
  );


  and

  (
    g373_p,
    a_1__p_spl_01,
    b_4__p_spl_11
  );


  or

  (
    g373_n,
    a_1__n_spl_01,
    b_4__n_spl_11
  );


  and

  (
    g374_p,
    g325_p_spl_0,
    g373_p_spl_0
  );


  or

  (
    g374_n,
    g325_n_spl_0,
    g373_n_spl_0
  );


  and

  (
    g375_p,
    g325_n_spl_,
    g373_n_spl_0
  );


  or

  (
    g375_n,
    g325_p_spl_,
    g373_p_spl_0
  );


  and

  (
    g376_p,
    g374_n_spl_,
    g375_n
  );


  or

  (
    g376_n,
    g374_p_spl_,
    g375_p
  );


  and

  (
    g377_p,
    g372_p_spl_,
    g376_p_spl_
  );


  or

  (
    g377_n,
    g372_n_spl_,
    g376_n_spl_
  );


  and

  (
    g378_p,
    g372_n_spl_,
    g376_n_spl_
  );


  or

  (
    g378_n,
    g372_p_spl_,
    g376_p_spl_
  );


  and

  (
    g379_p,
    g377_n_spl_,
    g378_n
  );


  or

  (
    g379_n,
    g377_p_spl_,
    g378_p
  );


  and

  (
    g380_p,
    g368_p_spl_,
    g370_n_spl_
  );


  or

  (
    g380_n,
    g368_n_spl_,
    g370_p_spl_
  );


  and

  (
    g381_p,
    g371_n_spl_,
    g380_n
  );


  or

  (
    g381_n,
    g371_p_spl_,
    g380_p
  );


  and

  (
    g382_p,
    g379_p_spl_,
    g381_p_spl_
  );


  or

  (
    g382_n,
    g379_n_spl_,
    g381_n_spl_
  );


  and

  (
    g383_p,
    g371_n_spl_,
    g382_n_spl_
  );


  or

  (
    g383_n,
    g371_p_spl_,
    g382_p_spl_
  );


  and

  (
    g384_p,
    g333_n_spl_,
    g335_n_spl_
  );


  or

  (
    g384_n,
    g333_p_spl_,
    g335_p_spl_
  );


  and

  (
    g385_p,
    g336_n_spl_,
    g384_n
  );


  or

  (
    g385_n,
    g336_p_spl_,
    g384_p
  );


  and

  (
    g386_p,
    g383_n_spl_,
    g385_p_spl_
  );


  or

  (
    g386_n,
    g383_p_spl_,
    g385_n_spl_
  );


  and

  (
    g387_p,
    g374_n_spl_,
    g377_n_spl_
  );


  or

  (
    g387_n,
    g374_p_spl_,
    g377_p_spl_
  );


  and

  (
    g388_p,
    a_0__p_spl_01,
    b_6__p_spl_11
  );


  or

  (
    g388_n,
    a_0__n_spl_01,
    b_6__n_spl_11
  );


  and

  (
    g389_p,
    g387_n_spl_,
    g388_p_spl_
  );


  or

  (
    g389_n,
    g387_p_spl_,
    g388_n_spl_
  );


  and

  (
    g390_p,
    g387_p_spl_,
    g388_n_spl_
  );


  or

  (
    g390_n,
    g387_n_spl_,
    g388_p_spl_
  );


  and

  (
    g391_p,
    g389_n_spl_0,
    g390_n
  );


  or

  (
    g391_n,
    g389_p_spl_0,
    g390_p
  );


  and

  (
    g392_p,
    g383_p_spl_,
    g385_n_spl_
  );


  or

  (
    g392_n,
    g383_n_spl_,
    g385_p_spl_
  );


  and

  (
    g393_p,
    g386_n_spl_,
    g392_n
  );


  or

  (
    g393_n,
    g386_p_spl_,
    g392_p
  );


  and

  (
    g394_p,
    g391_p_spl_,
    g393_p_spl_
  );


  or

  (
    g394_n,
    g391_n_spl_,
    g393_n_spl_
  );


  and

  (
    g395_p,
    g386_n_spl_,
    g394_n_spl_
  );


  or

  (
    g395_n,
    g386_p_spl_,
    g394_p_spl_
  );


  and

  (
    g396_p,
    g346_n_spl_,
    g348_n_spl_
  );


  or

  (
    g396_n,
    g346_p_spl_,
    g348_p_spl_
  );


  and

  (
    g397_p,
    g349_n_spl_,
    g396_n
  );


  or

  (
    g397_n,
    g349_p_spl_,
    g396_p
  );


  and

  (
    g398_p,
    g395_n_spl_,
    g397_p_spl_
  );


  or

  (
    g398_n,
    g395_p_spl_,
    g397_n_spl_
  );


  and

  (
    g399_p,
    g395_p_spl_,
    g397_n_spl_
  );


  or

  (
    g399_n,
    g395_n_spl_,
    g397_p_spl_
  );


  and

  (
    g400_p,
    g398_n_spl_,
    g399_n
  );


  or

  (
    g400_n,
    g398_p_spl_,
    g399_p
  );


  and

  (
    g401_p,
    g389_p_spl_0,
    g400_p_spl_
  );


  or

  (
    g401_n,
    g389_n_spl_0,
    g400_n_spl_
  );


  and

  (
    g402_p,
    g398_n_spl_,
    g401_n_spl_
  );


  or

  (
    g402_n,
    g398_p_spl_,
    g401_p_spl_
  );


  and

  (
    g403_p,
    g344_n_spl_,
    g355_n_spl_
  );


  or

  (
    g403_n,
    g344_p_spl_,
    g355_p_spl_
  );


  and

  (
    g404_p,
    g356_n_spl_,
    g403_n
  );


  or

  (
    g404_n,
    g356_p_spl_,
    g403_p
  );


  and

  (
    g405_p,
    g402_n_spl_,
    g404_p_spl_
  );


  or

  (
    g405_n,
    g402_p_spl_,
    g404_n_spl_
  );


  and

  (
    g406_p,
    a_2__p_spl_11,
    b_0__p_spl_10
  );


  or

  (
    g406_n,
    a_2__n_spl_11,
    b_0__n_spl_10
  );


  and

  (
    g407_p,
    g362_p_spl_,
    g406_p_spl_0
  );


  or

  (
    g407_n,
    g362_n_spl_,
    g406_n_spl_0
  );


  and

  (
    g408_p,
    a_1__p_spl_10,
    b_2__p_spl_11
  );


  or

  (
    g408_n,
    a_1__n_spl_10,
    b_2__n_spl_11
  );


  and

  (
    g409_p,
    a_3__p_spl_11,
    b_0__p_spl_10
  );


  or

  (
    g409_n,
    a_3__n_spl_11,
    b_0__n_spl_11
  );


  and

  (
    g410_p,
    a_2__p_spl_11,
    b_1__p_spl_10
  );


  or

  (
    g410_n,
    a_2__n_spl_11,
    b_1__n_spl_11
  );


  and

  (
    g411_p,
    g409_n,
    g410_n
  );


  or

  (
    g411_n,
    g409_p,
    g410_p
  );


  and

  (
    g412_p,
    g407_n_spl_,
    g411_n
  );


  or

  (
    g412_n,
    g407_p_spl_,
    g411_p
  );


  and

  (
    g413_p,
    g408_p_spl_,
    g412_p_spl_
  );


  or

  (
    g413_n,
    g408_n_spl_,
    g412_n_spl_
  );


  and

  (
    g414_p,
    g407_n_spl_,
    g413_n_spl_
  );


  or

  (
    g414_n,
    g407_p_spl_,
    g413_p_spl_
  );


  and

  (
    g415_p,
    g364_n_spl_,
    g366_n_spl_
  );


  or

  (
    g415_n,
    g364_p_spl_,
    g366_p_spl_
  );


  and

  (
    g416_p,
    g367_n_spl_,
    g415_n
  );


  or

  (
    g416_n,
    g367_p_spl_,
    g415_p
  );


  and

  (
    g417_p,
    g414_n_spl_,
    g416_p_spl_
  );


  or

  (
    g417_n,
    g414_p_spl_,
    g416_n_spl_
  );


  and

  (
    g418_p,
    a_0__p_spl_01,
    b_3__p_spl_11
  );


  or

  (
    g418_n,
    a_0__n_spl_01,
    b_3__n_spl_11
  );


  and

  (
    g419_p,
    g373_p_spl_,
    g418_p_spl_0
  );


  or

  (
    g419_n,
    g373_n_spl_,
    g418_n_spl_0
  );


  and

  (
    g420_p,
    a_1__p_spl_10,
    b_3__p_spl_11
  );


  or

  (
    g420_n,
    a_1__n_spl_10,
    b_3__n_spl_11
  );


  and

  (
    g421_p,
    a_0__p_spl_10,
    b_4__p_spl_11
  );


  or

  (
    g421_n,
    a_0__n_spl_10,
    b_4__n_spl_11
  );


  and

  (
    g422_p,
    g420_n,
    g421_n
  );


  or

  (
    g422_n,
    g420_p,
    g421_p
  );


  and

  (
    g423_p,
    g419_n_spl_0,
    g422_n
  );


  or

  (
    g423_n,
    g419_p_spl_0,
    g422_p
  );


  and

  (
    g424_p,
    g414_p_spl_,
    g416_n_spl_
  );


  or

  (
    g424_n,
    g414_n_spl_,
    g416_p_spl_
  );


  and

  (
    g425_p,
    g417_n_spl_,
    g424_n
  );


  or

  (
    g425_n,
    g417_p_spl_,
    g424_p
  );


  and

  (
    g426_p,
    g423_p_spl_,
    g425_p_spl_
  );


  or

  (
    g426_n,
    g423_n_spl_,
    g425_n_spl_
  );


  and

  (
    g427_p,
    g417_n_spl_,
    g426_n_spl_
  );


  or

  (
    g427_n,
    g417_p_spl_,
    g426_p_spl_
  );


  and

  (
    g428_p,
    g379_n_spl_,
    g381_n_spl_
  );


  or

  (
    g428_n,
    g379_p_spl_,
    g381_p_spl_
  );


  and

  (
    g429_p,
    g382_n_spl_,
    g428_n
  );


  or

  (
    g429_n,
    g382_p_spl_,
    g428_p
  );


  and

  (
    g430_p,
    g427_n_spl_,
    g429_p_spl_
  );


  or

  (
    g430_n,
    g427_p_spl_,
    g429_n_spl_
  );


  and

  (
    g431_p,
    g427_p_spl_,
    g429_n_spl_
  );


  or

  (
    g431_n,
    g427_n_spl_,
    g429_p_spl_
  );


  and

  (
    g432_p,
    g430_n_spl_,
    g431_n
  );


  or

  (
    g432_n,
    g430_p_spl_,
    g431_p
  );


  and

  (
    g433_p,
    g419_p_spl_0,
    g432_p_spl_
  );


  or

  (
    g433_n,
    g419_n_spl_0,
    g432_n_spl_
  );


  and

  (
    g434_p,
    g430_n_spl_,
    g433_n_spl_
  );


  or

  (
    g434_n,
    g430_p_spl_,
    g433_p_spl_
  );


  and

  (
    g435_p,
    g391_n_spl_,
    g393_n_spl_
  );


  or

  (
    g435_n,
    g391_p_spl_,
    g393_p_spl_
  );


  and

  (
    g436_p,
    g394_n_spl_,
    g435_n
  );


  or

  (
    g436_n,
    g394_p_spl_,
    g435_p
  );


  and

  (
    g437_p,
    g434_n_spl_,
    g436_p_spl_
  );


  or

  (
    g437_n,
    g434_p_spl_,
    g436_n_spl_
  );


  and

  (
    g438_p,
    g389_n_spl_,
    g400_n_spl_
  );


  or

  (
    g438_n,
    g389_p_spl_,
    g400_p_spl_
  );


  and

  (
    g439_p,
    g401_n_spl_,
    g438_n
  );


  or

  (
    g439_n,
    g401_p_spl_,
    g438_p
  );


  and

  (
    g440_p,
    g437_p_spl_0,
    g439_p_spl_
  );


  or

  (
    g440_n,
    g437_n_spl_0,
    g439_n_spl_
  );


  and

  (
    g441_p,
    g437_n_spl_0,
    g439_n_spl_
  );


  or

  (
    g441_n,
    g437_p_spl_0,
    g439_p_spl_
  );


  and

  (
    g442_p,
    g440_n_spl_,
    g441_n
  );


  or

  (
    g442_n,
    g440_p_spl_,
    g441_p
  );


  and

  (
    g443_p,
    g434_p_spl_,
    g436_n_spl_
  );


  or

  (
    g443_n,
    g434_n_spl_,
    g436_p_spl_
  );


  and

  (
    g444_p,
    g437_n_spl_,
    g443_n
  );


  or

  (
    g444_n,
    g437_p_spl_,
    g443_p
  );


  and

  (
    g445_p,
    a_1__p_spl_11,
    b_1__p_spl_11
  );


  or

  (
    g445_n,
    a_1__n_spl_1,
    b_1__n_spl_11
  );


  and

  (
    g446_p,
    g406_p_spl_0,
    g445_p_spl_0
  );


  or

  (
    g446_n,
    g406_n_spl_0,
    g445_n_spl_0
  );


  and

  (
    g447_p,
    a_0__p_spl_10,
    b_2__p_spl_11
  );


  or

  (
    g447_n,
    a_0__n_spl_10,
    b_2__n_spl_11
  );


  and

  (
    g448_p,
    g406_n_spl_,
    g445_n_spl_0
  );


  or

  (
    g448_n,
    g406_p_spl_,
    g445_p_spl_0
  );


  and

  (
    g449_p,
    g446_n_spl_,
    g448_n
  );


  or

  (
    g449_n,
    g446_p_spl_,
    g448_p
  );


  and

  (
    g450_p,
    g447_p_spl_,
    g449_p_spl_
  );


  or

  (
    g450_n,
    g447_n_spl_,
    g449_n_spl_
  );


  and

  (
    g451_p,
    g446_n_spl_,
    g450_n_spl_
  );


  or

  (
    g451_n,
    g446_p_spl_,
    g450_p_spl_
  );


  and

  (
    g452_p,
    g408_n_spl_,
    g412_n_spl_
  );


  or

  (
    g452_n,
    g408_p_spl_,
    g412_p_spl_
  );


  and

  (
    g453_p,
    g413_n_spl_,
    g452_n
  );


  or

  (
    g453_n,
    g413_p_spl_,
    g452_p
  );


  and

  (
    g454_p,
    g451_n_spl_,
    g453_p_spl_
  );


  or

  (
    g454_n,
    g451_p_spl_,
    g453_n_spl_
  );


  and

  (
    g455_p,
    g451_p_spl_,
    g453_n_spl_
  );


  or

  (
    g455_n,
    g451_n_spl_,
    g453_p_spl_
  );


  and

  (
    g456_p,
    g454_n_spl_,
    g455_n
  );


  or

  (
    g456_n,
    g454_p_spl_,
    g455_p
  );


  and

  (
    g457_p,
    g418_p_spl_0,
    g456_p_spl_
  );


  or

  (
    g457_n,
    g418_n_spl_0,
    g456_n_spl_
  );


  and

  (
    g458_p,
    g454_n_spl_,
    g457_n_spl_
  );


  or

  (
    g458_n,
    g454_p_spl_,
    g457_p_spl_
  );


  and

  (
    g459_p,
    g423_n_spl_,
    g425_n_spl_
  );


  or

  (
    g459_n,
    g423_p_spl_,
    g425_p_spl_
  );


  and

  (
    g460_p,
    g426_n_spl_,
    g459_n
  );


  or

  (
    g460_n,
    g426_p_spl_,
    g459_p
  );


  and

  (
    g461_p,
    g458_n_spl_,
    g460_p_spl_
  );


  or

  (
    g461_n,
    g458_p_spl_,
    g460_n_spl_
  );


  and

  (
    g462_p,
    g419_n_spl_,
    g432_n_spl_
  );


  or

  (
    g462_n,
    g419_p_spl_,
    g432_p_spl_
  );


  and

  (
    g463_p,
    g433_n_spl_,
    g462_n
  );


  or

  (
    g463_n,
    g433_p_spl_,
    g462_p
  );


  and

  (
    g464_p,
    g461_p_spl_0,
    g463_p_spl_0
  );


  or

  (
    g464_n,
    g461_n_spl_0,
    g463_n_spl_0
  );


  and

  (
    g465_p,
    a_0__p_spl_11,
    b_0__p_spl_11
  );


  or

  (
    g465_n,
    a_0__n_spl_1,
    b_0__n_spl_11
  );


  and

  (
    g466_p,
    g445_p_spl_,
    g465_p_spl_
  );


  or

  (
    g466_n,
    g445_n_spl_,
    g465_n
  );


  and

  (
    g467_p,
    g447_n_spl_,
    g449_n_spl_
  );


  or

  (
    g467_n,
    g447_p_spl_,
    g449_p_spl_
  );


  and

  (
    g468_p,
    g450_n_spl_,
    g467_n
  );


  or

  (
    g468_n,
    g450_p_spl_,
    g467_p
  );


  and

  (
    g469_p,
    g466_p_spl_,
    g468_p_spl_
  );


  or

  (
    g469_n,
    g466_n_spl_,
    g468_n
  );


  and

  (
    g470_p,
    g418_n_spl_,
    g456_n_spl_
  );


  or

  (
    g470_n,
    g418_p_spl_,
    g456_p_spl_
  );


  and

  (
    g471_p,
    g457_n_spl_,
    g470_n
  );


  or

  (
    g471_n,
    g457_p_spl_,
    g470_p
  );


  and

  (
    g472_p,
    g469_p_spl_,
    g471_p_spl_
  );


  or

  (
    g472_n,
    g469_n_spl_,
    g471_n
  );


  and

  (
    g473_p,
    g458_p_spl_,
    g460_n_spl_
  );


  or

  (
    g473_n,
    g458_n_spl_,
    g460_p_spl_
  );


  and

  (
    g474_p,
    g461_n_spl_0,
    g473_n
  );


  or

  (
    g474_n,
    g461_p_spl_0,
    g473_p
  );


  and

  (
    g475_p,
    g472_p_spl_,
    g474_p_spl_
  );


  or

  (
    g475_n,
    g472_n_spl_,
    g474_n
  );


  and

  (
    g476_p,
    g463_p_spl_0,
    g475_p_spl_
  );


  or

  (
    g476_n,
    g463_n_spl_0,
    g475_n_spl_0
  );


  and

  (
    g477_p,
    g464_n,
    g476_n
  );


  or

  (
    g477_n,
    g464_p,
    g476_p
  );


  and

  (
    g478_p,
    g444_p_spl_,
    g477_n_spl_
  );


  or

  (
    g478_n,
    g444_n,
    g477_p
  );


  and

  (
    g479_p,
    g442_p_spl_,
    g478_p_spl_
  );


  or

  (
    g479_n,
    g442_n,
    g478_n_spl_
  );


  and

  (
    g480_p,
    g440_n_spl_,
    g479_n_spl_
  );


  or

  (
    g480_n,
    g440_p_spl_,
    g479_p
  );


  and

  (
    g481_p,
    g402_p_spl_,
    g404_n_spl_
  );


  or

  (
    g481_n,
    g402_n_spl_,
    g404_p_spl_
  );


  and

  (
    g482_p,
    g405_n_spl_,
    g481_n
  );


  or

  (
    g482_n,
    g405_p_spl_,
    g481_p
  );


  and

  (
    g483_p,
    g480_n_spl_,
    g482_p_spl_
  );


  or

  (
    g483_n,
    g480_p,
    g482_n
  );


  and

  (
    g484_p,
    g405_n_spl_,
    g483_n_spl_
  );


  or

  (
    g484_n,
    g405_p_spl_,
    g483_p
  );


  and

  (
    g485_p,
    g357_p_spl_,
    g359_n_spl_
  );


  or

  (
    g485_n,
    g357_n_spl_,
    g359_p_spl_
  );


  and

  (
    g486_p,
    g360_n_spl_,
    g485_n
  );


  or

  (
    g486_n,
    g360_p_spl_,
    g485_p
  );


  and

  (
    g487_p,
    g484_n_spl_,
    g486_p_spl_
  );


  or

  (
    g487_n,
    g484_p,
    g486_n
  );


  and

  (
    g488_p,
    g360_n_spl_,
    g487_n_spl_
  );


  or

  (
    g488_n,
    g360_p_spl_,
    g487_p
  );


  and

  (
    g489_p,
    g314_p_spl_,
    g488_n_spl_
  );


  or

  (
    g489_n,
    g314_n,
    g488_p
  );


  and

  (
    g490_p,
    g312_n_spl_,
    g489_n_spl_
  );


  or

  (
    g490_n,
    g312_p_spl_,
    g489_p
  );


  and

  (
    g491_p,
    g251_p_spl_,
    g490_n_spl_
  );


  or

  (
    g491_n,
    g251_n,
    g490_p
  );


  and

  (
    g492_p,
    g249_n_spl_,
    g491_n_spl_
  );


  or

  (
    g492_n,
    g249_p_spl_,
    g491_p
  );


  and

  (
    g493_p,
    g193_p_spl_,
    g195_n_spl_
  );


  or

  (
    g493_n,
    g193_n_spl_,
    g195_p_spl_
  );


  and

  (
    g494_p,
    g196_n_spl_,
    g493_n
  );


  or

  (
    g494_n,
    g196_p_spl_,
    g493_p
  );


  and

  (
    g495_p,
    g492_n_spl_,
    g494_p_spl_
  );


  or

  (
    g495_n,
    g492_p,
    g494_n
  );


  and

  (
    g496_p,
    g196_n_spl_,
    g495_n_spl_
  );


  or

  (
    g496_n,
    g196_p_spl_,
    g495_p
  );


  and

  (
    g497_p,
    g149_n_spl_,
    g496_n_spl_
  );


  or

  (
    g497_n,
    g149_p_spl_,
    g496_p_spl_
  );


  and

  (
    g498_p,
    g148_n_spl_,
    g497_n
  );


  or

  (
    g498_n,
    g148_p_spl_,
    g497_p
  );


  and

  (
    g499_p,
    g107_p_spl_,
    g498_n_spl_
  );


  or

  (
    g499_n,
    g107_n,
    g498_p
  );


  or

  (
    g500_n,
    g30_p_spl_,
    g48_p_spl_
  );


  or

  (
    g501_n,
    g99_p_spl_,
    g102_p_spl_
  );


  and

  (
    g502_p,
    g500_n,
    g501_n
  );


  or

  (
    g503_n,
    g105_p_spl_,
    g502_p
  );


  or

  (
    g504_n,
    g499_p,
    g503_n
  );


  or

  (
    g505_n,
    g49_p,
    g504_n
  );


  and

  (
    g506_p,
    g148_n_spl_,
    g149_n_spl_
  );


  or

  (
    g506_n,
    g148_p_spl_,
    g149_p_spl_
  );


  and

  (
    g507_p,
    g496_n_spl_,
    g506_n
  );


  and

  (
    g508_p,
    g496_p_spl_,
    g506_p
  );


  or

  (
    g509_n,
    g507_p,
    g508_p
  );


  or

  (
    g510_n,
    g492_n_spl_,
    g494_p_spl_
  );


  and

  (
    g511_p,
    g495_n_spl_,
    g510_n
  );


  or

  (
    g512_n,
    g251_p_spl_,
    g490_n_spl_
  );


  and

  (
    g513_p,
    g491_n_spl_,
    g512_n
  );


  and

  (
    g514_p,
    g511_p_spl_,
    g513_p_spl_
  );


  or

  (
    g515_n,
    g314_p_spl_,
    g488_n_spl_
  );


  and

  (
    g516_p,
    g489_n_spl_,
    g515_n
  );


  or

  (
    g517_n,
    g484_n_spl_,
    g486_p_spl_
  );


  and

  (
    g518_p,
    g487_n_spl_,
    g517_n
  );


  or

  (
    g519_n,
    g480_n_spl_,
    g482_p_spl_
  );


  and

  (
    g520_p,
    g483_n_spl_,
    g519_n
  );


  or

  (
    g521_n,
    g442_p_spl_,
    g478_p_spl_
  );


  and

  (
    g522_p,
    g479_n_spl_,
    g521_n
  );


  and

  (
    g523_p,
    g520_p_spl_,
    g522_p_spl_
  );


  and

  (
    g524_p,
    g518_p_spl_,
    g523_p
  );


  and

  (
    g525_p,
    g516_p_spl_,
    g524_p
  );


  and

  (
    g526_p,
    g514_p,
    g525_p
  );


  and

  (
    g527_p,
    g509_n_spl_,
    g526_p
  );


  or

  (
    g528_n,
    g505_n_spl_0,
    g527_p
  );


  or

  (
    g529_n,
    g107_p_spl_,
    g498_n_spl_
  );


  and

  (
    g530_p,
    g499_n,
    g529_n
  );


  or

  (
    g531_n,
    g513_p_spl_,
    g516_p_spl_
  );


  or

  (
    g532_n,
    g518_p_spl_,
    g520_p_spl_
  );


  or

  (
    g533_n,
    g522_p_spl_,
    g532_n
  );


  or

  (
    g534_n,
    g511_p_spl_,
    g533_n
  );


  or

  (
    g535_n,
    g509_n_spl_,
    g534_n
  );


  or

  (
    g536_n,
    g531_n,
    g535_n
  );


  or

  (
    g537_n,
    g530_p,
    g536_n
  );


  and

  (
    g538_p,
    g505_n_spl_0,
    g537_n
  );


  or

  (
    g539_n,
    g465_p_spl_,
    g538_p_spl_00
  );


  and

  (
    g540_p,
    g528_n_spl_00,
    g539_n
  );


  and

  (
    g541_p,
    a_1__p_spl_11,
    b_0__p_spl_11
  );


  and

  (
    g542_p,
    a_0__p_spl_11,
    b_1__p_spl_11
  );


  or

  (
    g543_n,
    g541_p,
    g542_p
  );


  and

  (
    g544_p,
    g466_n_spl_,
    g543_n
  );


  and

  (
    g545_p,
    g528_n_spl_00,
    g544_p
  );


  or

  (
    g546_n,
    g538_p_spl_00,
    g545_p
  );


  or

  (
    g547_n,
    g466_p_spl_,
    g468_p_spl_
  );


  and

  (
    g548_p,
    g469_n_spl_,
    g547_n
  );


  and

  (
    g549_p,
    g528_n_spl_01,
    g548_p
  );


  or

  (
    g550_n,
    g538_p_spl_01,
    g549_p
  );


  or

  (
    g551_n,
    g469_p_spl_,
    g471_p_spl_
  );


  and

  (
    g552_p,
    g472_n_spl_,
    g551_n
  );


  and

  (
    g553_p,
    g528_n_spl_01,
    g552_p
  );


  or

  (
    g554_n,
    g538_p_spl_01,
    g553_p
  );


  or

  (
    g555_n,
    g472_p_spl_,
    g474_p_spl_
  );


  and

  (
    g556_p,
    g475_n_spl_0,
    g555_n
  );


  and

  (
    g557_p,
    g528_n_spl_10,
    g556_p
  );


  or

  (
    g558_n,
    g538_p_spl_10,
    g557_p
  );


  and

  (
    g559_p,
    g461_n_spl_,
    g475_n_spl_
  );


  or

  (
    g559_n,
    g461_p_spl_,
    g475_p_spl_
  );


  and

  (
    g560_p,
    g463_p_spl_,
    g559_p
  );


  and

  (
    g561_p,
    g463_n_spl_,
    g559_n
  );


  or

  (
    g562_n,
    g560_p,
    g561_p
  );


  and

  (
    g563_p,
    g528_n_spl_10,
    g562_n
  );


  or

  (
    g564_n,
    g538_p_spl_10,
    g563_p
  );


  or

  (
    g565_n,
    g444_p_spl_,
    g477_n_spl_
  );


  and

  (
    g566_p,
    g478_n_spl_,
    g565_n
  );


  and

  (
    g567_p,
    g528_n_spl_1,
    g566_p
  );


  or

  (
    g568_n,
    g538_p_spl_1,
    g567_p
  );


  buf

  (
    product_0_,
    g540_p
  );


  buf

  (
    product_1_,
    g546_n
  );


  buf

  (
    product_2_,
    g550_n
  );


  buf

  (
    product_3_,
    g554_n
  );


  buf

  (
    product_4_,
    g558_n
  );


  buf

  (
    product_5_,
    g564_n
  );


  buf

  (
    product_6_,
    g568_n
  );


  not

  (
    product_7_,
    g505_n_spl_
  );


  buf

  (
    a_7__p_spl_,
    a_7__p
  );


  buf

  (
    a_7__p_spl_0,
    a_7__p_spl_
  );


  buf

  (
    a_7__p_spl_00,
    a_7__p_spl_0
  );


  buf

  (
    a_7__p_spl_01,
    a_7__p_spl_0
  );


  buf

  (
    a_7__p_spl_1,
    a_7__p_spl_
  );


  buf

  (
    a_7__p_spl_10,
    a_7__p_spl_1
  );


  buf

  (
    a_7__p_spl_11,
    a_7__p_spl_1
  );


  buf

  (
    b_4__p_spl_,
    b_4__p
  );


  buf

  (
    b_4__p_spl_0,
    b_4__p_spl_
  );


  buf

  (
    b_4__p_spl_00,
    b_4__p_spl_0
  );


  buf

  (
    b_4__p_spl_01,
    b_4__p_spl_0
  );


  buf

  (
    b_4__p_spl_1,
    b_4__p_spl_
  );


  buf

  (
    b_4__p_spl_10,
    b_4__p_spl_1
  );


  buf

  (
    b_4__p_spl_11,
    b_4__p_spl_1
  );


  buf

  (
    a_7__n_spl_,
    a_7__n
  );


  buf

  (
    a_7__n_spl_0,
    a_7__n_spl_
  );


  buf

  (
    a_7__n_spl_00,
    a_7__n_spl_0
  );


  buf

  (
    a_7__n_spl_01,
    a_7__n_spl_0
  );


  buf

  (
    a_7__n_spl_1,
    a_7__n_spl_
  );


  buf

  (
    a_7__n_spl_10,
    a_7__n_spl_1
  );


  buf

  (
    a_7__n_spl_11,
    a_7__n_spl_1
  );


  buf

  (
    b_4__n_spl_,
    b_4__n
  );


  buf

  (
    b_4__n_spl_0,
    b_4__n_spl_
  );


  buf

  (
    b_4__n_spl_00,
    b_4__n_spl_0
  );


  buf

  (
    b_4__n_spl_01,
    b_4__n_spl_0
  );


  buf

  (
    b_4__n_spl_1,
    b_4__n_spl_
  );


  buf

  (
    b_4__n_spl_10,
    b_4__n_spl_1
  );


  buf

  (
    b_4__n_spl_11,
    b_4__n_spl_1
  );


  buf

  (
    b_3__p_spl_,
    b_3__p
  );


  buf

  (
    b_3__p_spl_0,
    b_3__p_spl_
  );


  buf

  (
    b_3__p_spl_00,
    b_3__p_spl_0
  );


  buf

  (
    b_3__p_spl_000,
    b_3__p_spl_00
  );


  buf

  (
    b_3__p_spl_01,
    b_3__p_spl_0
  );


  buf

  (
    b_3__p_spl_1,
    b_3__p_spl_
  );


  buf

  (
    b_3__p_spl_10,
    b_3__p_spl_1
  );


  buf

  (
    b_3__p_spl_11,
    b_3__p_spl_1
  );


  buf

  (
    g17_p_spl_,
    g17_p
  );


  buf

  (
    g17_p_spl_0,
    g17_p_spl_
  );


  buf

  (
    b_3__n_spl_,
    b_3__n
  );


  buf

  (
    b_3__n_spl_0,
    b_3__n_spl_
  );


  buf

  (
    b_3__n_spl_00,
    b_3__n_spl_0
  );


  buf

  (
    b_3__n_spl_000,
    b_3__n_spl_00
  );


  buf

  (
    b_3__n_spl_01,
    b_3__n_spl_0
  );


  buf

  (
    b_3__n_spl_1,
    b_3__n_spl_
  );


  buf

  (
    b_3__n_spl_10,
    b_3__n_spl_1
  );


  buf

  (
    b_3__n_spl_11,
    b_3__n_spl_1
  );


  buf

  (
    g17_n_spl_,
    g17_n
  );


  buf

  (
    g17_n_spl_0,
    g17_n_spl_
  );


  buf

  (
    g19_n_spl_,
    g19_n
  );


  buf

  (
    g19_p_spl_,
    g19_p
  );


  buf

  (
    g18_n_spl_,
    g18_n
  );


  buf

  (
    g18_n_spl_0,
    g18_n_spl_
  );


  buf

  (
    g18_p_spl_,
    g18_p
  );


  buf

  (
    g18_p_spl_0,
    g18_p_spl_
  );


  buf

  (
    b_5__p_spl_,
    b_5__p
  );


  buf

  (
    b_5__p_spl_0,
    b_5__p_spl_
  );


  buf

  (
    b_5__p_spl_00,
    b_5__p_spl_0
  );


  buf

  (
    b_5__p_spl_01,
    b_5__p_spl_0
  );


  buf

  (
    b_5__p_spl_1,
    b_5__p_spl_
  );


  buf

  (
    b_5__p_spl_10,
    b_5__p_spl_1
  );


  buf

  (
    b_5__p_spl_11,
    b_5__p_spl_1
  );


  buf

  (
    b_5__n_spl_,
    b_5__n
  );


  buf

  (
    b_5__n_spl_0,
    b_5__n_spl_
  );


  buf

  (
    b_5__n_spl_00,
    b_5__n_spl_0
  );


  buf

  (
    b_5__n_spl_01,
    b_5__n_spl_0
  );


  buf

  (
    b_5__n_spl_1,
    b_5__n_spl_
  );


  buf

  (
    b_5__n_spl_10,
    b_5__n_spl_1
  );


  buf

  (
    b_5__n_spl_11,
    b_5__n_spl_1
  );


  buf

  (
    g21_p_spl_,
    g21_p
  );


  buf

  (
    g21_p_spl_0,
    g21_p_spl_
  );


  buf

  (
    g21_p_spl_1,
    g21_p_spl_
  );


  buf

  (
    g22_p_spl_,
    g22_p
  );


  buf

  (
    g21_n_spl_,
    g21_n
  );


  buf

  (
    g21_n_spl_0,
    g21_n_spl_
  );


  buf

  (
    g21_n_spl_1,
    g21_n_spl_
  );


  buf

  (
    g22_n_spl_,
    g22_n
  );


  buf

  (
    g23_n_spl_,
    g23_n
  );


  buf

  (
    g23_p_spl_,
    g23_p
  );


  buf

  (
    b_6__p_spl_,
    b_6__p
  );


  buf

  (
    b_6__p_spl_0,
    b_6__p_spl_
  );


  buf

  (
    b_6__p_spl_00,
    b_6__p_spl_0
  );


  buf

  (
    b_6__p_spl_01,
    b_6__p_spl_0
  );


  buf

  (
    b_6__p_spl_1,
    b_6__p_spl_
  );


  buf

  (
    b_6__p_spl_10,
    b_6__p_spl_1
  );


  buf

  (
    b_6__p_spl_11,
    b_6__p_spl_1
  );


  buf

  (
    b_6__n_spl_,
    b_6__n
  );


  buf

  (
    b_6__n_spl_0,
    b_6__n_spl_
  );


  buf

  (
    b_6__n_spl_00,
    b_6__n_spl_0
  );


  buf

  (
    b_6__n_spl_01,
    b_6__n_spl_0
  );


  buf

  (
    b_6__n_spl_1,
    b_6__n_spl_
  );


  buf

  (
    b_6__n_spl_10,
    b_6__n_spl_1
  );


  buf

  (
    b_6__n_spl_11,
    b_6__n_spl_1
  );


  buf

  (
    a_6__n_spl_,
    a_6__n
  );


  buf

  (
    a_6__n_spl_0,
    a_6__n_spl_
  );


  buf

  (
    a_6__n_spl_00,
    a_6__n_spl_0
  );


  buf

  (
    a_6__n_spl_01,
    a_6__n_spl_0
  );


  buf

  (
    a_6__n_spl_1,
    a_6__n_spl_
  );


  buf

  (
    a_6__n_spl_10,
    a_6__n_spl_1
  );


  buf

  (
    a_6__n_spl_11,
    a_6__n_spl_1
  );


  buf

  (
    b_7__p_spl_,
    b_7__p
  );


  buf

  (
    b_7__p_spl_0,
    b_7__p_spl_
  );


  buf

  (
    b_7__p_spl_00,
    b_7__p_spl_0
  );


  buf

  (
    b_7__p_spl_000,
    b_7__p_spl_00
  );


  buf

  (
    b_7__p_spl_001,
    b_7__p_spl_00
  );


  buf

  (
    b_7__p_spl_01,
    b_7__p_spl_0
  );


  buf

  (
    b_7__p_spl_1,
    b_7__p_spl_
  );


  buf

  (
    b_7__p_spl_10,
    b_7__p_spl_1
  );


  buf

  (
    b_7__p_spl_11,
    b_7__p_spl_1
  );


  buf

  (
    a_6__p_spl_,
    a_6__p
  );


  buf

  (
    a_6__p_spl_0,
    a_6__p_spl_
  );


  buf

  (
    a_6__p_spl_00,
    a_6__p_spl_0
  );


  buf

  (
    a_6__p_spl_01,
    a_6__p_spl_0
  );


  buf

  (
    a_6__p_spl_1,
    a_6__p_spl_
  );


  buf

  (
    a_6__p_spl_10,
    a_6__p_spl_1
  );


  buf

  (
    a_6__p_spl_11,
    a_6__p_spl_1
  );


  buf

  (
    b_7__n_spl_,
    b_7__n
  );


  buf

  (
    b_7__n_spl_0,
    b_7__n_spl_
  );


  buf

  (
    b_7__n_spl_00,
    b_7__n_spl_0
  );


  buf

  (
    b_7__n_spl_000,
    b_7__n_spl_00
  );


  buf

  (
    b_7__n_spl_001,
    b_7__n_spl_00
  );


  buf

  (
    b_7__n_spl_01,
    b_7__n_spl_0
  );


  buf

  (
    b_7__n_spl_1,
    b_7__n_spl_
  );


  buf

  (
    b_7__n_spl_10,
    b_7__n_spl_1
  );


  buf

  (
    b_7__n_spl_11,
    b_7__n_spl_1
  );


  buf

  (
    g25_p_spl_,
    g25_p
  );


  buf

  (
    g26_n_spl_,
    g26_n
  );


  buf

  (
    g25_n_spl_,
    g25_n
  );


  buf

  (
    g26_p_spl_,
    g26_p
  );


  buf

  (
    g27_n_spl_,
    g27_n
  );


  buf

  (
    g27_p_spl_,
    g27_p
  );


  buf

  (
    g24_p_spl_,
    g24_p
  );


  buf

  (
    g24_p_spl_0,
    g24_p_spl_
  );


  buf

  (
    g24_p_spl_1,
    g24_p_spl_
  );


  buf

  (
    g29_p_spl_,
    g29_p
  );


  buf

  (
    g24_n_spl_,
    g24_n
  );


  buf

  (
    g24_n_spl_0,
    g24_n_spl_
  );


  buf

  (
    g24_n_spl_1,
    g24_n_spl_
  );


  buf

  (
    g29_n_spl_,
    g29_n
  );


  buf

  (
    b_0__p_spl_,
    b_0__p
  );


  buf

  (
    b_0__p_spl_0,
    b_0__p_spl_
  );


  buf

  (
    b_0__p_spl_00,
    b_0__p_spl_0
  );


  buf

  (
    b_0__p_spl_000,
    b_0__p_spl_00
  );


  buf

  (
    b_0__p_spl_01,
    b_0__p_spl_0
  );


  buf

  (
    b_0__p_spl_1,
    b_0__p_spl_
  );


  buf

  (
    b_0__p_spl_10,
    b_0__p_spl_1
  );


  buf

  (
    b_0__p_spl_11,
    b_0__p_spl_1
  );


  buf

  (
    b_0__n_spl_,
    b_0__n
  );


  buf

  (
    b_0__n_spl_0,
    b_0__n_spl_
  );


  buf

  (
    b_0__n_spl_00,
    b_0__n_spl_0
  );


  buf

  (
    b_0__n_spl_01,
    b_0__n_spl_0
  );


  buf

  (
    b_0__n_spl_1,
    b_0__n_spl_
  );


  buf

  (
    b_0__n_spl_10,
    b_0__n_spl_1
  );


  buf

  (
    b_0__n_spl_11,
    b_0__n_spl_1
  );


  buf

  (
    b_1__p_spl_,
    b_1__p
  );


  buf

  (
    b_1__p_spl_0,
    b_1__p_spl_
  );


  buf

  (
    b_1__p_spl_00,
    b_1__p_spl_0
  );


  buf

  (
    b_1__p_spl_000,
    b_1__p_spl_00
  );


  buf

  (
    b_1__p_spl_01,
    b_1__p_spl_0
  );


  buf

  (
    b_1__p_spl_1,
    b_1__p_spl_
  );


  buf

  (
    b_1__p_spl_10,
    b_1__p_spl_1
  );


  buf

  (
    b_1__p_spl_11,
    b_1__p_spl_1
  );


  buf

  (
    g33_p_spl_,
    g33_p
  );


  buf

  (
    g33_p_spl_0,
    g33_p_spl_
  );


  buf

  (
    b_1__n_spl_,
    b_1__n
  );


  buf

  (
    b_1__n_spl_0,
    b_1__n_spl_
  );


  buf

  (
    b_1__n_spl_00,
    b_1__n_spl_0
  );


  buf

  (
    b_1__n_spl_01,
    b_1__n_spl_0
  );


  buf

  (
    b_1__n_spl_1,
    b_1__n_spl_
  );


  buf

  (
    b_1__n_spl_10,
    b_1__n_spl_1
  );


  buf

  (
    b_1__n_spl_11,
    b_1__n_spl_1
  );


  buf

  (
    g33_n_spl_,
    g33_n
  );


  buf

  (
    g33_n_spl_0,
    g33_n_spl_
  );


  buf

  (
    b_2__p_spl_,
    b_2__p
  );


  buf

  (
    b_2__p_spl_0,
    b_2__p_spl_
  );


  buf

  (
    b_2__p_spl_00,
    b_2__p_spl_0
  );


  buf

  (
    b_2__p_spl_000,
    b_2__p_spl_00
  );


  buf

  (
    b_2__p_spl_01,
    b_2__p_spl_0
  );


  buf

  (
    b_2__p_spl_1,
    b_2__p_spl_
  );


  buf

  (
    b_2__p_spl_10,
    b_2__p_spl_1
  );


  buf

  (
    b_2__p_spl_11,
    b_2__p_spl_1
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g34_p_spl_0,
    g34_p_spl_
  );


  buf

  (
    b_2__n_spl_,
    b_2__n
  );


  buf

  (
    b_2__n_spl_0,
    b_2__n_spl_
  );


  buf

  (
    b_2__n_spl_00,
    b_2__n_spl_0
  );


  buf

  (
    b_2__n_spl_000,
    b_2__n_spl_00
  );


  buf

  (
    b_2__n_spl_01,
    b_2__n_spl_0
  );


  buf

  (
    b_2__n_spl_1,
    b_2__n_spl_
  );


  buf

  (
    b_2__n_spl_10,
    b_2__n_spl_1
  );


  buf

  (
    b_2__n_spl_11,
    b_2__n_spl_1
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g34_n_spl_0,
    g34_n_spl_
  );


  buf

  (
    g32_p_spl_,
    g32_p
  );


  buf

  (
    g32_p_spl_0,
    g32_p_spl_
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    g35_p_spl_0,
    g35_p_spl_
  );


  buf

  (
    g35_p_spl_00,
    g35_p_spl_0
  );


  buf

  (
    g35_p_spl_01,
    g35_p_spl_0
  );


  buf

  (
    g35_p_spl_1,
    g35_p_spl_
  );


  buf

  (
    g35_p_spl_10,
    g35_p_spl_1
  );


  buf

  (
    g32_n_spl_,
    g32_n
  );


  buf

  (
    g32_n_spl_0,
    g32_n_spl_
  );


  buf

  (
    g35_n_spl_,
    g35_n
  );


  buf

  (
    g35_n_spl_0,
    g35_n_spl_
  );


  buf

  (
    g35_n_spl_00,
    g35_n_spl_0
  );


  buf

  (
    g35_n_spl_01,
    g35_n_spl_0
  );


  buf

  (
    g35_n_spl_1,
    g35_n_spl_
  );


  buf

  (
    g35_n_spl_10,
    g35_n_spl_1
  );


  buf

  (
    g37_n_spl_,
    g37_n
  );


  buf

  (
    g39_n_spl_,
    g39_n
  );


  buf

  (
    g39_n_spl_0,
    g39_n_spl_
  );


  buf

  (
    g37_p_spl_,
    g37_p
  );


  buf

  (
    g39_p_spl_,
    g39_p
  );


  buf

  (
    g39_p_spl_0,
    g39_p_spl_
  );


  buf

  (
    g40_n_spl_,
    g40_n
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g41_n_spl_,
    g41_n
  );


  buf

  (
    g41_n_spl_0,
    g41_n_spl_
  );


  buf

  (
    g41_n_spl_00,
    g41_n_spl_0
  );


  buf

  (
    g41_n_spl_01,
    g41_n_spl_0
  );


  buf

  (
    g41_n_spl_1,
    g41_n_spl_
  );


  buf

  (
    g41_p_spl_,
    g41_p
  );


  buf

  (
    g41_p_spl_0,
    g41_p_spl_
  );


  buf

  (
    g41_p_spl_00,
    g41_p_spl_0
  );


  buf

  (
    g41_p_spl_01,
    g41_p_spl_0
  );


  buf

  (
    g41_p_spl_1,
    g41_p_spl_
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    g36_n_spl_,
    g36_n
  );


  buf

  (
    g36_n_spl_0,
    g36_n_spl_
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g30_p_spl_,
    g30_p
  );


  buf

  (
    g30_p_spl_0,
    g30_p_spl_
  );


  buf

  (
    g44_p_spl_,
    g44_p
  );


  buf

  (
    g44_p_spl_0,
    g44_p_spl_
  );


  buf

  (
    g44_p_spl_1,
    g44_p_spl_
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    g44_n_spl_,
    g44_n
  );


  buf

  (
    g44_n_spl_0,
    g44_n_spl_
  );


  buf

  (
    g44_n_spl_1,
    g44_n_spl_
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    g48_p_spl_,
    g48_p
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    g52_n_spl_,
    g52_n
  );


  buf

  (
    g53_n_spl_,
    g53_n
  );


  buf

  (
    g53_p_spl_,
    g53_p
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g56_n_spl_,
    g56_n
  );


  buf

  (
    g56_p_spl_,
    g56_p
  );


  buf

  (
    g51_p_spl_,
    g51_p
  );


  buf

  (
    g57_n_spl_,
    g57_n
  );


  buf

  (
    g51_n_spl_,
    g51_n
  );


  buf

  (
    g57_p_spl_,
    g57_p
  );


  buf

  (
    a_5__p_spl_,
    a_5__p
  );


  buf

  (
    a_5__p_spl_0,
    a_5__p_spl_
  );


  buf

  (
    a_5__p_spl_00,
    a_5__p_spl_0
  );


  buf

  (
    a_5__p_spl_01,
    a_5__p_spl_0
  );


  buf

  (
    a_5__p_spl_1,
    a_5__p_spl_
  );


  buf

  (
    a_5__p_spl_10,
    a_5__p_spl_1
  );


  buf

  (
    a_5__p_spl_11,
    a_5__p_spl_1
  );


  buf

  (
    a_5__n_spl_,
    a_5__n
  );


  buf

  (
    a_5__n_spl_0,
    a_5__n_spl_
  );


  buf

  (
    a_5__n_spl_00,
    a_5__n_spl_0
  );


  buf

  (
    a_5__n_spl_01,
    a_5__n_spl_0
  );


  buf

  (
    a_5__n_spl_1,
    a_5__n_spl_
  );


  buf

  (
    a_5__n_spl_10,
    a_5__n_spl_1
  );


  buf

  (
    a_5__n_spl_11,
    a_5__n_spl_1
  );


  buf

  (
    a_4__n_spl_,
    a_4__n
  );


  buf

  (
    a_4__n_spl_0,
    a_4__n_spl_
  );


  buf

  (
    a_4__n_spl_00,
    a_4__n_spl_0
  );


  buf

  (
    a_4__n_spl_01,
    a_4__n_spl_0
  );


  buf

  (
    a_4__n_spl_1,
    a_4__n_spl_
  );


  buf

  (
    a_4__n_spl_10,
    a_4__n_spl_1
  );


  buf

  (
    a_4__n_spl_11,
    a_4__n_spl_1
  );


  buf

  (
    a_4__p_spl_,
    a_4__p
  );


  buf

  (
    a_4__p_spl_0,
    a_4__p_spl_
  );


  buf

  (
    a_4__p_spl_00,
    a_4__p_spl_0
  );


  buf

  (
    a_4__p_spl_01,
    a_4__p_spl_0
  );


  buf

  (
    a_4__p_spl_1,
    a_4__p_spl_
  );


  buf

  (
    a_4__p_spl_10,
    a_4__p_spl_1
  );


  buf

  (
    a_4__p_spl_11,
    a_4__p_spl_1
  );


  buf

  (
    g59_p_spl_,
    g59_p
  );


  buf

  (
    g60_p_spl_,
    g60_p
  );


  buf

  (
    g59_n_spl_,
    g59_n
  );


  buf

  (
    g60_n_spl_,
    g60_n
  );


  buf

  (
    g63_p_spl_,
    g63_p
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g63_n_spl_,
    g63_n
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    g65_n_spl_0,
    g65_n_spl_
  );


  buf

  (
    g65_p_spl_,
    g65_p
  );


  buf

  (
    g65_p_spl_0,
    g65_p_spl_
  );


  buf

  (
    g62_n_spl_,
    g62_n
  );


  buf

  (
    g67_p_spl_,
    g67_p
  );


  buf

  (
    g62_p_spl_,
    g62_p
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    g68_n_spl_,
    g68_n
  );


  buf

  (
    g68_p_spl_,
    g68_p
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g61_p_spl_0,
    g61_p_spl_
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g61_n_spl_0,
    g61_n_spl_
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    g71_n_spl_,
    g71_n
  );


  buf

  (
    g71_p_spl_,
    g71_p
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    g79_p_spl_,
    g79_p
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    g82_p_spl_,
    g82_p
  );


  buf

  (
    g82_n_spl_,
    g82_n
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g83_p_spl_,
    g83_p
  );


  buf

  (
    g85_p_spl_,
    g85_p
  );


  buf

  (
    g85_n_spl_,
    g85_n
  );


  buf

  (
    g86_n_spl_,
    g86_n
  );


  buf

  (
    g86_p_spl_,
    g86_p
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    g89_n_spl_,
    g89_n
  );


  buf

  (
    g89_p_spl_,
    g89_p
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g93_n_spl_,
    g93_n
  );


  buf

  (
    g93_p_spl_,
    g93_p
  );


  buf

  (
    g97_n_spl_,
    g97_n
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    g97_p_spl_,
    g97_p
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    g99_p_spl_,
    g99_p
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    g101_p_spl_,
    g101_p
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g101_n_spl_,
    g101_n
  );


  buf

  (
    g102_p_spl_,
    g102_p
  );


  buf

  (
    g94_n_spl_,
    g94_n
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g94_p_spl_,
    g94_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g105_p_spl_,
    g105_p
  );


  buf

  (
    g109_p_spl_,
    g109_p
  );


  buf

  (
    g109_n_spl_,
    g109_n
  );


  buf

  (
    g111_n_spl_,
    g111_n
  );


  buf

  (
    g111_p_spl_,
    g111_p
  );


  buf

  (
    g110_n_spl_,
    g110_n
  );


  buf

  (
    g110_p_spl_,
    g110_p
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    g113_p_spl_,
    g113_p
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    g113_n_spl_,
    g113_n
  );


  buf

  (
    g114_n_spl_,
    g114_n
  );


  buf

  (
    g114_p_spl_,
    g114_p
  );


  buf

  (
    g116_p_spl_,
    g116_p
  );


  buf

  (
    g116_n_spl_,
    g116_n
  );


  buf

  (
    g117_n_spl_,
    g117_n
  );


  buf

  (
    g117_p_spl_,
    g117_p
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g120_p_spl_,
    g120_p
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g120_n_spl_,
    g120_n
  );


  buf

  (
    a_3__n_spl_,
    a_3__n
  );


  buf

  (
    a_3__n_spl_0,
    a_3__n_spl_
  );


  buf

  (
    a_3__n_spl_00,
    a_3__n_spl_0
  );


  buf

  (
    a_3__n_spl_01,
    a_3__n_spl_0
  );


  buf

  (
    a_3__n_spl_1,
    a_3__n_spl_
  );


  buf

  (
    a_3__n_spl_10,
    a_3__n_spl_1
  );


  buf

  (
    a_3__n_spl_11,
    a_3__n_spl_1
  );


  buf

  (
    a_3__p_spl_,
    a_3__p
  );


  buf

  (
    a_3__p_spl_0,
    a_3__p_spl_
  );


  buf

  (
    a_3__p_spl_00,
    a_3__p_spl_0
  );


  buf

  (
    a_3__p_spl_01,
    a_3__p_spl_0
  );


  buf

  (
    a_3__p_spl_1,
    a_3__p_spl_
  );


  buf

  (
    a_3__p_spl_10,
    a_3__p_spl_1
  );


  buf

  (
    a_3__p_spl_11,
    a_3__p_spl_1
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g123_p_spl_,
    g123_p
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    g123_n_spl_,
    g123_n
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    g128_n_spl_,
    g128_n
  );


  buf

  (
    g128_p_spl_,
    g128_p
  );


  buf

  (
    g124_p_spl_,
    g124_p
  );


  buf

  (
    g124_p_spl_0,
    g124_p_spl_
  );


  buf

  (
    g130_p_spl_,
    g130_p
  );


  buf

  (
    g124_n_spl_,
    g124_n
  );


  buf

  (
    g124_n_spl_0,
    g124_n_spl_
  );


  buf

  (
    g130_n_spl_,
    g130_n
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g135_p_spl_,
    g135_p
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g135_n_spl_,
    g135_n
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g136_p_spl_,
    g136_p
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    g139_p_spl_,
    g139_p
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    g139_n_spl_,
    g139_n
  );


  buf

  (
    g140_n_spl_,
    g140_n
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g141_n_spl_,
    g141_n
  );


  buf

  (
    g143_p_spl_,
    g143_p
  );


  buf

  (
    g141_p_spl_,
    g141_p
  );


  buf

  (
    g143_n_spl_,
    g143_n
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g145_n_spl_,
    g145_n
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g145_p_spl_,
    g145_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g151_p_spl_,
    g151_p
  );


  buf

  (
    g151_p_spl_0,
    g151_p_spl_
  );


  buf

  (
    g151_p_spl_1,
    g151_p_spl_
  );


  buf

  (
    g151_n_spl_,
    g151_n
  );


  buf

  (
    g151_n_spl_0,
    g151_n_spl_
  );


  buf

  (
    g151_n_spl_1,
    g151_n_spl_
  );


  buf

  (
    g152_n_spl_,
    g152_n
  );


  buf

  (
    g152_p_spl_,
    g152_p
  );


  buf

  (
    g150_p_spl_,
    g150_p
  );


  buf

  (
    g155_p_spl_,
    g155_p
  );


  buf

  (
    g150_n_spl_,
    g150_n
  );


  buf

  (
    g155_n_spl_,
    g155_n
  );


  buf

  (
    g156_n_spl_,
    g156_n
  );


  buf

  (
    g156_p_spl_,
    g156_p
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g159_n_spl_0,
    g159_n_spl_
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g159_p_spl_0,
    g159_p_spl_
  );


  buf

  (
    g158_p_spl_,
    g158_p
  );


  buf

  (
    g164_p_spl_,
    g164_p
  );


  buf

  (
    g158_n_spl_,
    g158_n
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g166_n_spl_,
    g166_n
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g166_p_spl_,
    g166_p
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    a_2__n_spl_,
    a_2__n
  );


  buf

  (
    a_2__n_spl_0,
    a_2__n_spl_
  );


  buf

  (
    a_2__n_spl_00,
    a_2__n_spl_0
  );


  buf

  (
    a_2__n_spl_01,
    a_2__n_spl_0
  );


  buf

  (
    a_2__n_spl_1,
    a_2__n_spl_
  );


  buf

  (
    a_2__n_spl_10,
    a_2__n_spl_1
  );


  buf

  (
    a_2__n_spl_11,
    a_2__n_spl_1
  );


  buf

  (
    a_2__p_spl_,
    a_2__p
  );


  buf

  (
    a_2__p_spl_0,
    a_2__p_spl_
  );


  buf

  (
    a_2__p_spl_00,
    a_2__p_spl_0
  );


  buf

  (
    a_2__p_spl_01,
    a_2__p_spl_0
  );


  buf

  (
    a_2__p_spl_1,
    a_2__p_spl_
  );


  buf

  (
    a_2__p_spl_10,
    a_2__p_spl_1
  );


  buf

  (
    a_2__p_spl_11,
    a_2__p_spl_1
  );


  buf

  (
    g170_p_spl_,
    g170_p
  );


  buf

  (
    g171_p_spl_,
    g171_p
  );


  buf

  (
    g170_n_spl_,
    g170_n
  );


  buf

  (
    g171_n_spl_,
    g171_n
  );


  buf

  (
    g173_n_spl_,
    g173_n
  );


  buf

  (
    g175_p_spl_,
    g175_p
  );


  buf

  (
    g173_p_spl_,
    g173_p
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g176_n_spl_,
    g176_n
  );


  buf

  (
    g176_p_spl_,
    g176_p
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g172_p_spl_0,
    g172_p_spl_
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g172_n_spl_0,
    g172_n_spl_
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g179_p_spl_,
    g179_p
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g183_p_spl_,
    g183_p
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g183_n_spl_,
    g183_n
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g184_p_spl_,
    g184_p
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g188_n_spl_,
    g188_n
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g189_n_spl_,
    g189_n
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g189_p_spl_,
    g189_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g192_n_spl_,
    g192_n
  );


  buf

  (
    g192_p_spl_,
    g192_p
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g195_n_spl_,
    g195_n
  );


  buf

  (
    g197_n_spl_,
    g197_n
  );


  buf

  (
    g197_p_spl_,
    g197_p
  );


  buf

  (
    g198_p_spl_,
    g198_p
  );


  buf

  (
    g198_p_spl_0,
    g198_p_spl_
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    g198_n_spl_,
    g198_n
  );


  buf

  (
    g198_n_spl_0,
    g198_n_spl_
  );


  buf

  (
    g200_n_spl_,
    g200_n
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g203_p_spl_,
    g203_p
  );


  buf

  (
    g203_n_spl_,
    g203_n
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g209_p_spl_,
    g209_p
  );


  buf

  (
    g209_n_spl_,
    g209_n
  );


  buf

  (
    g210_n_spl_,
    g210_n
  );


  buf

  (
    g210_p_spl_,
    g210_p
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g212_p_spl_,
    g212_p
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g212_n_spl_,
    g212_n
  );


  buf

  (
    g213_n_spl_,
    g213_n
  );


  buf

  (
    g213_p_spl_,
    g213_p
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g215_p_spl_,
    g215_p
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g215_n_spl_,
    g215_n
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g218_n_spl_,
    g218_n
  );


  buf

  (
    g218_p_spl_,
    g218_p
  );


  buf

  (
    g219_n_spl_,
    g219_n
  );


  buf

  (
    g221_p_spl_,
    g221_p
  );


  buf

  (
    g219_p_spl_,
    g219_p
  );


  buf

  (
    g221_n_spl_,
    g221_n
  );


  buf

  (
    a_1__n_spl_,
    a_1__n
  );


  buf

  (
    a_1__n_spl_0,
    a_1__n_spl_
  );


  buf

  (
    a_1__n_spl_00,
    a_1__n_spl_0
  );


  buf

  (
    a_1__n_spl_01,
    a_1__n_spl_0
  );


  buf

  (
    a_1__n_spl_1,
    a_1__n_spl_
  );


  buf

  (
    a_1__n_spl_10,
    a_1__n_spl_1
  );


  buf

  (
    a_1__p_spl_,
    a_1__p
  );


  buf

  (
    a_1__p_spl_0,
    a_1__p_spl_
  );


  buf

  (
    a_1__p_spl_00,
    a_1__p_spl_0
  );


  buf

  (
    a_1__p_spl_01,
    a_1__p_spl_0
  );


  buf

  (
    a_1__p_spl_1,
    a_1__p_spl_
  );


  buf

  (
    a_1__p_spl_10,
    a_1__p_spl_1
  );


  buf

  (
    a_1__p_spl_11,
    a_1__p_spl_1
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g223_p_spl_0,
    g223_p_spl_
  );


  buf

  (
    g224_p_spl_,
    g224_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g223_n_spl_0,
    g223_n_spl_
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    g228_p_spl_,
    g228_p
  );


  buf

  (
    g226_p_spl_,
    g226_p
  );


  buf

  (
    g228_n_spl_,
    g228_n
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g225_p_spl_,
    g225_p
  );


  buf

  (
    g225_p_spl_0,
    g225_p_spl_
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g225_n_spl_,
    g225_n
  );


  buf

  (
    g225_n_spl_0,
    g225_n_spl_
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g232_n_spl_,
    g232_n
  );


  buf

  (
    g232_p_spl_,
    g232_p
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    g222_p_spl_,
    g222_p
  );


  buf

  (
    g234_p_spl_,
    g234_p
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g234_n_spl_,
    g234_n
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g237_n_spl_,
    g237_n
  );


  buf

  (
    g237_p_spl_,
    g237_p
  );


  buf

  (
    g238_n_spl_,
    g238_n
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    g241_p_spl_,
    g241_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g244_n_spl_,
    g244_n
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g246_n_spl_,
    g246_n
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g246_p_spl_,
    g246_p
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g249_n_spl_,
    g249_n
  );


  buf

  (
    g249_p_spl_,
    g249_p
  );


  buf

  (
    g252_p_spl_,
    g252_p
  );


  buf

  (
    g252_p_spl_0,
    g252_p_spl_
  );


  buf

  (
    g252_n_spl_,
    g252_n
  );


  buf

  (
    g252_n_spl_0,
    g252_n_spl_
  );


  buf

  (
    g253_n_spl_,
    g253_n
  );


  buf

  (
    g253_p_spl_,
    g253_p
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g254_p_spl_0,
    g254_p_spl_
  );


  buf

  (
    g258_p_spl_,
    g258_p
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g254_n_spl_0,
    g254_n_spl_
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g262_p_spl_,
    g262_p
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g262_n_spl_,
    g262_n
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g264_p_spl_,
    g264_p
  );


  buf

  (
    g264_p_spl_0,
    g264_p_spl_
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g264_n_spl_,
    g264_n
  );


  buf

  (
    g264_n_spl_0,
    g264_n_spl_
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g270_n_spl_,
    g270_n
  );


  buf

  (
    g270_p_spl_,
    g270_p
  );


  buf

  (
    g263_n_spl_,
    g263_n
  );


  buf

  (
    g263_p_spl_,
    g263_p
  );


  buf

  (
    g272_p_spl_,
    g272_p
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_p_spl_,
    g275_p
  );


  buf

  (
    g276_n_spl_,
    g276_n
  );


  buf

  (
    g278_p_spl_,
    g278_p
  );


  buf

  (
    g276_p_spl_,
    g276_p
  );


  buf

  (
    g278_n_spl_,
    g278_n
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g280_p_spl_0,
    g280_p_spl_
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g280_n_spl_0,
    g280_n_spl_
  );


  buf

  (
    a_0__n_spl_,
    a_0__n
  );


  buf

  (
    a_0__n_spl_0,
    a_0__n_spl_
  );


  buf

  (
    a_0__n_spl_00,
    a_0__n_spl_0
  );


  buf

  (
    a_0__n_spl_01,
    a_0__n_spl_0
  );


  buf

  (
    a_0__n_spl_1,
    a_0__n_spl_
  );


  buf

  (
    a_0__n_spl_10,
    a_0__n_spl_1
  );


  buf

  (
    a_0__p_spl_,
    a_0__p
  );


  buf

  (
    a_0__p_spl_0,
    a_0__p_spl_
  );


  buf

  (
    a_0__p_spl_00,
    a_0__p_spl_0
  );


  buf

  (
    a_0__p_spl_01,
    a_0__p_spl_0
  );


  buf

  (
    a_0__p_spl_1,
    a_0__p_spl_
  );


  buf

  (
    a_0__p_spl_10,
    a_0__p_spl_1
  );


  buf

  (
    a_0__p_spl_11,
    a_0__p_spl_1
  );


  buf

  (
    g281_n_spl_,
    g281_n
  );


  buf

  (
    g281_p_spl_,
    g281_p
  );


  buf

  (
    g282_p_spl_,
    g282_p
  );


  buf

  (
    g286_p_spl_,
    g286_p
  );


  buf

  (
    g282_n_spl_,
    g282_n
  );


  buf

  (
    g286_n_spl_,
    g286_n
  );


  buf

  (
    g287_n_spl_,
    g287_n
  );


  buf

  (
    g287_p_spl_,
    g287_p
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g291_p_spl_,
    g291_p
  );


  buf

  (
    g289_p_spl_,
    g289_p
  );


  buf

  (
    g291_n_spl_,
    g291_n
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g288_n_spl_,
    g288_n
  );


  buf

  (
    g294_p_spl_,
    g294_p
  );


  buf

  (
    g288_p_spl_,
    g288_p
  );


  buf

  (
    g294_n_spl_,
    g294_n
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g295_p_spl_,
    g295_p
  );


  buf

  (
    g279_n_spl_,
    g279_n
  );


  buf

  (
    g279_p_spl_,
    g279_p
  );


  buf

  (
    g297_p_spl_,
    g297_p
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g297_n_spl_,
    g297_n
  );


  buf

  (
    g299_n_spl_,
    g299_n
  );


  buf

  (
    g300_n_spl_,
    g300_n
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g301_p_spl_,
    g301_p
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g304_n_spl_,
    g304_n
  );


  buf

  (
    g304_p_spl_,
    g304_p
  );


  buf

  (
    g305_n_spl_,
    g305_n
  );


  buf

  (
    g307_p_spl_,
    g307_p
  );


  buf

  (
    g305_p_spl_,
    g305_p
  );


  buf

  (
    g307_n_spl_,
    g307_n
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    g308_p_spl_,
    g308_p
  );


  buf

  (
    g309_n_spl_,
    g309_n
  );


  buf

  (
    g311_p_spl_,
    g311_p
  );


  buf

  (
    g309_p_spl_,
    g309_p
  );


  buf

  (
    g311_n_spl_,
    g311_n
  );


  buf

  (
    g312_n_spl_,
    g312_n
  );


  buf

  (
    g312_p_spl_,
    g312_p
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g316_n_spl_,
    g316_n
  );


  buf

  (
    g316_p_spl_,
    g316_p
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g319_p_spl_,
    g319_p
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g319_n_spl_,
    g319_n
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g321_n_spl_,
    g321_n
  );


  buf

  (
    g323_p_spl_,
    g323_p
  );


  buf

  (
    g321_p_spl_,
    g321_p
  );


  buf

  (
    g323_n_spl_,
    g323_n
  );


  buf

  (
    g325_p_spl_,
    g325_p
  );


  buf

  (
    g325_p_spl_0,
    g325_p_spl_
  );


  buf

  (
    g325_n_spl_,
    g325_n
  );


  buf

  (
    g325_n_spl_0,
    g325_n_spl_
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    g326_p_spl_,
    g326_p
  );


  buf

  (
    g330_p_spl_,
    g330_p
  );


  buf

  (
    g330_n_spl_,
    g330_n
  );


  buf

  (
    g331_n_spl_,
    g331_n
  );


  buf

  (
    g331_p_spl_,
    g331_p
  );


  buf

  (
    g324_n_spl_,
    g324_n
  );


  buf

  (
    g324_p_spl_,
    g324_p
  );


  buf

  (
    g333_p_spl_,
    g333_p
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g333_n_spl_,
    g333_n
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g336_n_spl_,
    g336_n
  );


  buf

  (
    g336_p_spl_,
    g336_p
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g339_p_spl_,
    g339_p
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g339_n_spl_,
    g339_n
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g343_p_spl_,
    g343_p
  );


  buf

  (
    g341_p_spl_,
    g341_p
  );


  buf

  (
    g343_n_spl_,
    g343_n
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g344_n_spl_0,
    g344_n_spl_
  );


  buf

  (
    g344_p_spl_,
    g344_p
  );


  buf

  (
    g344_p_spl_0,
    g344_p_spl_
  );


  buf

  (
    g340_n_spl_,
    g340_n
  );


  buf

  (
    g340_p_spl_,
    g340_p
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g348_p_spl_,
    g348_p
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g348_n_spl_,
    g348_n
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g350_n_spl_,
    g350_n
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    g350_p_spl_,
    g350_p
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g353_n_spl_,
    g353_n
  );


  buf

  (
    g353_p_spl_,
    g353_p
  );


  buf

  (
    g355_p_spl_,
    g355_p
  );


  buf

  (
    g355_n_spl_,
    g355_n
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g356_p_spl_,
    g356_p
  );


  buf

  (
    g357_n_spl_,
    g357_n
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g357_p_spl_,
    g357_p
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g362_p_spl_,
    g362_p
  );


  buf

  (
    g362_p_spl_0,
    g362_p_spl_
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g362_n_spl_,
    g362_n
  );


  buf

  (
    g362_n_spl_0,
    g362_n_spl_
  );


  buf

  (
    g363_n_spl_,
    g363_n
  );


  buf

  (
    g363_p_spl_,
    g363_p
  );


  buf

  (
    g364_p_spl_,
    g364_p
  );


  buf

  (
    g366_p_spl_,
    g366_p
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    g366_n_spl_,
    g366_n
  );


  buf

  (
    g367_n_spl_,
    g367_n
  );


  buf

  (
    g367_p_spl_,
    g367_p
  );


  buf

  (
    g368_n_spl_,
    g368_n
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g368_p_spl_,
    g368_p
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g373_p_spl_0,
    g373_p_spl_
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g373_n_spl_0,
    g373_n_spl_
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    g377_p_spl_,
    g377_p
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    g371_p_spl_,
    g371_p
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g383_p_spl_,
    g383_p
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g389_n_spl_0,
    g389_n_spl_
  );


  buf

  (
    g389_p_spl_,
    g389_p
  );


  buf

  (
    g389_p_spl_0,
    g389_p_spl_
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g391_n_spl_,
    g391_n
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g394_p_spl_,
    g394_p
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g395_p_spl_,
    g395_p
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g398_n_spl_,
    g398_n
  );


  buf

  (
    g398_p_spl_,
    g398_p
  );


  buf

  (
    g400_p_spl_,
    g400_p
  );


  buf

  (
    g400_n_spl_,
    g400_n
  );


  buf

  (
    g401_n_spl_,
    g401_n
  );


  buf

  (
    g401_p_spl_,
    g401_p
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g404_p_spl_,
    g404_p
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g404_n_spl_,
    g404_n
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g406_p_spl_0,
    g406_p_spl_
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g407_n_spl_,
    g407_n
  );


  buf

  (
    g407_p_spl_,
    g407_p
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    g413_p_spl_,
    g413_p
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g418_p_spl_,
    g418_p
  );


  buf

  (
    g418_p_spl_0,
    g418_p_spl_
  );


  buf

  (
    g418_n_spl_,
    g418_n
  );


  buf

  (
    g418_n_spl_0,
    g418_n_spl_
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g419_n_spl_0,
    g419_n_spl_
  );


  buf

  (
    g419_p_spl_,
    g419_p
  );


  buf

  (
    g419_p_spl_0,
    g419_p_spl_
  );


  buf

  (
    g417_n_spl_,
    g417_n
  );


  buf

  (
    g417_p_spl_,
    g417_p
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g425_p_spl_,
    g425_p
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g425_n_spl_,
    g425_n
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g432_n_spl_,
    g432_n
  );


  buf

  (
    g433_n_spl_,
    g433_n
  );


  buf

  (
    g433_p_spl_,
    g433_p
  );


  buf

  (
    g434_n_spl_,
    g434_n
  );


  buf

  (
    g436_p_spl_,
    g436_p
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    g436_n_spl_,
    g436_n
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g437_p_spl_0,
    g437_p_spl_
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g437_n_spl_,
    g437_n
  );


  buf

  (
    g437_n_spl_0,
    g437_n_spl_
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g445_p_spl_,
    g445_p
  );


  buf

  (
    g445_p_spl_0,
    g445_p_spl_
  );


  buf

  (
    g445_n_spl_,
    g445_n
  );


  buf

  (
    g445_n_spl_0,
    g445_n_spl_
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g457_p_spl_,
    g457_p
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g460_n_spl_,
    g460_n
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g461_p_spl_0,
    g461_p_spl_
  );


  buf

  (
    g463_p_spl_,
    g463_p
  );


  buf

  (
    g463_p_spl_0,
    g463_p_spl_
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g461_n_spl_0,
    g461_n_spl_
  );


  buf

  (
    g463_n_spl_,
    g463_n
  );


  buf

  (
    g463_n_spl_0,
    g463_n_spl_
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g466_p_spl_,
    g466_p
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g466_n_spl_,
    g466_n
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g471_p_spl_,
    g471_p
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g474_p_spl_,
    g474_p
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g475_p_spl_,
    g475_p
  );


  buf

  (
    g475_n_spl_,
    g475_n
  );


  buf

  (
    g475_n_spl_0,
    g475_n_spl_
  );


  buf

  (
    g444_p_spl_,
    g444_p
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g483_n_spl_,
    g483_n
  );


  buf

  (
    g360_n_spl_,
    g360_n
  );


  buf

  (
    g360_p_spl_,
    g360_p
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g486_p_spl_,
    g486_p
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g314_p_spl_,
    g314_p
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g489_n_spl_,
    g489_n
  );


  buf

  (
    g251_p_spl_,
    g251_p
  );


  buf

  (
    g490_n_spl_,
    g490_n
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g492_n_spl_,
    g492_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g495_n_spl_,
    g495_n
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g496_n_spl_,
    g496_n
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g496_p_spl_,
    g496_p
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g107_p_spl_,
    g107_p
  );


  buf

  (
    g498_n_spl_,
    g498_n
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g520_p_spl_,
    g520_p
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g516_p_spl_,
    g516_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g505_n_spl_0,
    g505_n_spl_
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g538_p_spl_0,
    g538_p_spl_
  );


  buf

  (
    g538_p_spl_00,
    g538_p_spl_0
  );


  buf

  (
    g538_p_spl_01,
    g538_p_spl_0
  );


  buf

  (
    g538_p_spl_1,
    g538_p_spl_
  );


  buf

  (
    g538_p_spl_10,
    g538_p_spl_1
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g528_n_spl_0,
    g528_n_spl_
  );


  buf

  (
    g528_n_spl_00,
    g528_n_spl_0
  );


  buf

  (
    g528_n_spl_01,
    g528_n_spl_0
  );


  buf

  (
    g528_n_spl_1,
    g528_n_spl_
  );


  buf

  (
    g528_n_spl_10,
    g528_n_spl_1
  );


endmodule
