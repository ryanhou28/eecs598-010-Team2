module c499(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,
  G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,
  G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,G481,G482,
  G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,
  G498,G499,G5,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41;
output G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,G481,
  G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,
  G497,G498,G499;

  wire G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,
    G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,
    G175,G176,G177,G178,G179,G180,G181,G182,G183,G184,G185,G186,G189,G192,G195,
    G198,G201,G204,G207,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
    G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G247,
    G260,G273,G286,G299,G312,G325,G338,G339,G340,G341,G342,G343,G344,G345,G346,
    G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,G361,
    G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,
    G377,G378,G379,G380,G381,G382,G383,G384,G385,G386,G391,G396,G401,G406,G411,
    G416,G421,G426,G431,G436,G437,G438,G439,G440,G441,G442,G443,G444,G445,G446,
    G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,G461,
    G462,G463,G464,G465,G466,G467;

  xor (G146,G1,G2);
  xor (G147,G3,G4);
  xor (G148,G5,G6);
  xor (G149,G7,G8);
  xor (G150,G9,G10);
  xor (G151,G11,G12);
  xor (G152,G13,G14);
  xor (G153,G15,G16);
  xor (G154,G17,G18);
  xor (G155,G19,G20);
  xor (G156,G21,G22);
  xor (G157,G23,G24);
  xor (G158,G25,G26);
  xor (G159,G27,G28);
  xor (G160,G29,G30);
  xor (G161,G31,G32);
  and (G162,G33,G41);
  and (G163,G34,G41);
  and (G164,G35,G41);
  and (G165,G36,G41);
  and (G166,G37,G41);
  and (G167,G38,G41);
  and (G168,G39,G41);
  and (G169,G40,G41);
  xor (G170,G1,G5);
  xor (G171,G9,G13);
  xor (G172,G2,G6);
  xor (G173,G10,G14);
  xor (G174,G3,G7);
  xor (G175,G11,G15);
  xor (G176,G4,G8);
  xor (G177,G12,G16);
  xor (G178,G17,G21);
  xor (G179,G25,G29);
  xor (G180,G18,G22);
  xor (G181,G26,G30);
  xor (G182,G19,G23);
  xor (G183,G27,G31);
  xor (G184,G20,G24);
  xor (G185,G28,G32);
  xor (G186,G146,G147);
  xor (G189,G148,G149);
  xor (G192,G150,G151);
  xor (G195,G152,G153);
  xor (G198,G154,G155);
  xor (G201,G156,G157);
  xor (G204,G158,G159);
  xor (G207,G160,G161);
  xor (G210,G170,G171);
  xor (G211,G172,G173);
  xor (G212,G174,G175);
  xor (G213,G176,G177);
  xor (G214,G178,G179);
  xor (G215,G180,G181);
  xor (G216,G182,G183);
  xor (G217,G184,G185);
  xor (G218,G186,G189);
  xor (G219,G192,G195);
  xor (G220,G186,G192);
  xor (G221,G189,G195);
  xor (G222,G198,G201);
  xor (G223,G204,G207);
  xor (G224,G198,G204);
  xor (G225,G201,G207);
  xor (G226,G162,G222);
  xor (G227,G163,G223);
  xor (G228,G164,G224);
  xor (G229,G165,G225);
  xor (G230,G166,G218);
  xor (G231,G167,G219);
  xor (G232,G168,G220);
  xor (G233,G169,G221);
  xor (G234,G210,G226);
  xor (G247,G211,G227);
  xor (G260,G212,G228);
  xor (G273,G213,G229);
  xor (G286,G214,G230);
  xor (G299,G215,G231);
  xor (G312,G216,G232);
  xor (G325,G217,G233);
  not (G338,G234);
  not (G339,G247);
  not (G340,G260);
  not (G341,G234);
  not (G342,G247);
  not (G343,G273);
  not (G344,G234);
  not (G345,G260);
  not (G346,G273);
  not (G347,G247);
  not (G348,G260);
  not (G349,G273);
  not (G350,G299);
  not (G351,G325);
  not (G352,G299);
  not (G353,G312);
  not (G354,G286);
  not (G355,G325);
  not (G356,G286);
  not (G357,G312);
  not (G358,G286);
  not (G359,G299);
  not (G360,G312);
  not (G361,G286);
  not (G362,G299);
  not (G363,G325);
  not (G364,G286);
  not (G365,G312);
  not (G366,G325);
  not (G367,G299);
  not (G368,G312);
  not (G369,G325);
  not (G370,G247);
  not (G371,G273);
  not (G372,G247);
  not (G373,G260);
  not (G374,G234);
  not (G375,G273);
  not (G376,G234);
  not (G377,G260);
  and (G378,G338,G339,G340,G273);
  and (G379,G341,G342,G260,G343);
  and (G380,G344,G247,G345,G346);
  and (G381,G234,G347,G348,G349);
  and (G382,G358,G359,G360,G325);
  and (G383,G361,G362,G312,G363);
  and (G384,G364,G299,G365,G366);
  and (G385,G286,G367,G368,G369);
  or (G386,G378,G379,G380,G381);
  or (G391,G382,G383,G384,G385);
  and (G396,G286,G350,G312,G351,G386);
  and (G401,G286,G352,G353,G325,G386);
  and (G406,G354,G299,G312,G355,G386);
  and (G411,G356,G299,G357,G325,G386);
  and (G416,G234,G370,G260,G371,G391);
  and (G421,G234,G372,G373,G273,G391);
  and (G426,G374,G247,G260,G375,G391);
  and (G431,G376,G247,G377,G273,G391);
  and (G436,G234,G396);
  and (G437,G247,G396);
  and (G438,G260,G396);
  and (G439,G273,G396);
  and (G440,G234,G401);
  and (G441,G247,G401);
  and (G442,G260,G401);
  and (G443,G273,G401);
  and (G444,G234,G406);
  and (G445,G247,G406);
  and (G446,G260,G406);
  and (G447,G273,G406);
  and (G448,G234,G411);
  and (G449,G247,G411);
  and (G450,G260,G411);
  and (G451,G273,G411);
  and (G452,G286,G416);
  and (G453,G299,G416);
  and (G454,G312,G416);
  and (G455,G325,G416);
  and (G456,G286,G421);
  and (G457,G299,G421);
  and (G458,G312,G421);
  and (G459,G325,G421);
  and (G460,G286,G426);
  and (G461,G299,G426);
  and (G462,G312,G426);
  and (G463,G325,G426);
  and (G464,G286,G431);
  and (G465,G299,G431);
  and (G466,G312,G431);
  and (G467,G325,G431);
  xor (G468,G1,G436);
  xor (G469,G2,G437);
  xor (G470,G3,G438);
  xor (G471,G4,G439);
  xor (G472,G5,G440);
  xor (G473,G6,G441);
  xor (G474,G7,G442);
  xor (G475,G8,G443);
  xor (G476,G9,G444);
  xor (G477,G10,G445);
  xor (G478,G11,G446);
  xor (G479,G12,G447);
  xor (G480,G13,G448);
  xor (G481,G14,G449);
  xor (G482,G15,G450);
  xor (G483,G16,G451);
  xor (G484,G17,G452);
  xor (G485,G18,G453);
  xor (G486,G19,G454);
  xor (G487,G20,G455);
  xor (G488,G21,G456);
  xor (G489,G22,G457);
  xor (G490,G23,G458);
  xor (G491,G24,G459);
  xor (G492,G25,G460);
  xor (G493,G26,G461);
  xor (G494,G27,G462);
  xor (G495,G28,G463);
  xor (G496,G29,G464);
  xor (G497,G30,G465);
  xor (G498,G31,G466);
  xor (G499,G32,G467);

endmodule
