
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  n630_lo,
  n642_lo,
  n654_lo,
  n666_lo,
  n678_lo,
  n690_lo,
  n702_lo,
  n714_lo,
  n726_lo,
  n738_lo,
  n750_lo,
  n762_lo,
  n774_lo,
  n786_lo,
  n798_lo,
  n810_lo,
  n822_lo,
  n834_lo,
  n846_lo,
  n858_lo,
  n870_lo,
  n882_lo,
  n894_lo,
  n906_lo,
  n918_lo,
  n930_lo,
  n942_lo,
  n954_lo,
  n966_lo,
  n978_lo,
  n990_lo,
  n1002_lo,
  n1005_lo,
  n1008_lo,
  n1017_lo,
  n1020_lo,
  n1029_lo,
  n1032_lo,
  n1041_lo,
  n1044_lo,
  n1053_lo,
  n1056_lo,
  n1065_lo,
  n1068_lo,
  n1077_lo,
  n1080_lo,
  n1089_lo,
  n1092_lo,
  n1101_lo,
  n1104_lo,
  n1837_o2,
  n1838_o2,
  n1839_o2,
  n1840_o2,
  n1841_o2,
  n1842_o2,
  n1843_o2,
  n1844_o2,
  n1845_o2,
  n1846_o2,
  n1847_o2,
  n1848_o2,
  n1849_o2,
  n1850_o2,
  n1851_o2,
  n1852_o2,
  n1853_o2,
  n1854_o2,
  n1855_o2,
  n1856_o2,
  n1857_o2,
  n1858_o2,
  n1859_o2,
  n1860_o2,
  n1861_o2,
  n1862_o2,
  n1863_o2,
  n1864_o2,
  n1865_o2,
  n1866_o2,
  n1867_o2,
  n1868_o2,
  G834_o2,
  G847_o2,
  G860_o2,
  G873_o2,
  G925_o2,
  G886_o2,
  G912_o2,
  G899_o2,
  n2151_o2,
  n2152_o2,
  n2153_o2,
  n2154_o2,
  n2155_o2,
  n2156_o2,
  n2157_o2,
  n2158_o2,
  n2159_o2,
  n2160_o2,
  n2161_o2,
  n2162_o2,
  n2163_o2,
  n2164_o2,
  n2165_o2,
  n2166_o2,
  n2167_o2,
  n2168_o2,
  n2169_o2,
  n2170_o2,
  n2171_o2,
  n2172_o2,
  n2173_o2,
  n2174_o2,
  n2175_o2,
  n2176_o2,
  n2177_o2,
  n2178_o2,
  n2179_o2,
  n2180_o2,
  n2181_o2,
  n2182_o2,
  G974_o2,
  G976_o2,
  G970_o2,
  G972_o2,
  G973_o2,
  G977_o2,
  G971_o2,
  G975_o2,
  G954_o2,
  G956_o2,
  G950_o2,
  G952_o2,
  G953_o2,
  G957_o2,
  G951_o2,
  G955_o2,
  G986_o2,
  G991_o2,
  G770_o2,
  G773_o2,
  G776_o2,
  G779_o2,
  G782_o2,
  G785_o2,
  G788_o2,
  G791_o2,
  G642_o2,
  G645_o2,
  G648_o2,
  G651_o2,
  G654_o2,
  G657_o2,
  G660_o2,
  G663_o2,
  G602_o2,
  G607_o2,
  G612_o2,
  G617_o2,
  G622_o2,
  G627_o2,
  G632_o2,
  G637_o2,
  n627_lo_buf_o2,
  n639_lo_buf_o2,
  n651_lo_buf_o2,
  n663_lo_buf_o2,
  n675_lo_buf_o2,
  n687_lo_buf_o2,
  n699_lo_buf_o2,
  n711_lo_buf_o2,
  n723_lo_buf_o2,
  n735_lo_buf_o2,
  n747_lo_buf_o2,
  n759_lo_buf_o2,
  n771_lo_buf_o2,
  n783_lo_buf_o2,
  n795_lo_buf_o2,
  n807_lo_buf_o2,
  n819_lo_buf_o2,
  n831_lo_buf_o2,
  n843_lo_buf_o2,
  n855_lo_buf_o2,
  n867_lo_buf_o2,
  n879_lo_buf_o2,
  n891_lo_buf_o2,
  n903_lo_buf_o2,
  n915_lo_buf_o2,
  n927_lo_buf_o2,
  n939_lo_buf_o2,
  n951_lo_buf_o2,
  n963_lo_buf_o2,
  n975_lo_buf_o2,
  n987_lo_buf_o2,
  n999_lo_buf_o2,
  G1324,
  G1325,
  G1326,
  G1327,
  G1328,
  G1329,
  G1330,
  G1331,
  G1332,
  G1333,
  G1334,
  G1335,
  G1336,
  G1337,
  G1338,
  G1339,
  G1340,
  G1341,
  G1342,
  G1343,
  G1344,
  G1345,
  G1346,
  G1347,
  G1348,
  G1349,
  G1350,
  G1351,
  G1352,
  G1353,
  G1354,
  G1355,
  n630_li,
  n642_li,
  n654_li,
  n666_li,
  n678_li,
  n690_li,
  n702_li,
  n714_li,
  n726_li,
  n738_li,
  n750_li,
  n762_li,
  n774_li,
  n786_li,
  n798_li,
  n810_li,
  n822_li,
  n834_li,
  n846_li,
  n858_li,
  n870_li,
  n882_li,
  n894_li,
  n906_li,
  n918_li,
  n930_li,
  n942_li,
  n954_li,
  n966_li,
  n978_li,
  n990_li,
  n1002_li,
  n1005_li,
  n1008_li,
  n1017_li,
  n1020_li,
  n1029_li,
  n1032_li,
  n1041_li,
  n1044_li,
  n1053_li,
  n1056_li,
  n1065_li,
  n1068_li,
  n1077_li,
  n1080_li,
  n1089_li,
  n1092_li,
  n1101_li,
  n1104_li,
  n1837_i2,
  n1838_i2,
  n1839_i2,
  n1840_i2,
  n1841_i2,
  n1842_i2,
  n1843_i2,
  n1844_i2,
  n1845_i2,
  n1846_i2,
  n1847_i2,
  n1848_i2,
  n1849_i2,
  n1850_i2,
  n1851_i2,
  n1852_i2,
  n1853_i2,
  n1854_i2,
  n1855_i2,
  n1856_i2,
  n1857_i2,
  n1858_i2,
  n1859_i2,
  n1860_i2,
  n1861_i2,
  n1862_i2,
  n1863_i2,
  n1864_i2,
  n1865_i2,
  n1866_i2,
  n1867_i2,
  n1868_i2,
  G834_i2,
  G847_i2,
  G860_i2,
  G873_i2,
  G925_i2,
  G886_i2,
  G912_i2,
  G899_i2,
  n2151_i2,
  n2152_i2,
  n2153_i2,
  n2154_i2,
  n2155_i2,
  n2156_i2,
  n2157_i2,
  n2158_i2,
  n2159_i2,
  n2160_i2,
  n2161_i2,
  n2162_i2,
  n2163_i2,
  n2164_i2,
  n2165_i2,
  n2166_i2,
  n2167_i2,
  n2168_i2,
  n2169_i2,
  n2170_i2,
  n2171_i2,
  n2172_i2,
  n2173_i2,
  n2174_i2,
  n2175_i2,
  n2176_i2,
  n2177_i2,
  n2178_i2,
  n2179_i2,
  n2180_i2,
  n2181_i2,
  n2182_i2,
  G974_i2,
  G976_i2,
  G970_i2,
  G972_i2,
  G973_i2,
  G977_i2,
  G971_i2,
  G975_i2,
  G954_i2,
  G956_i2,
  G950_i2,
  G952_i2,
  G953_i2,
  G957_i2,
  G951_i2,
  G955_i2,
  G986_i2,
  G991_i2,
  G770_i2,
  G773_i2,
  G776_i2,
  G779_i2,
  G782_i2,
  G785_i2,
  G788_i2,
  G791_i2,
  G642_i2,
  G645_i2,
  G648_i2,
  G651_i2,
  G654_i2,
  G657_i2,
  G660_i2,
  G663_i2,
  G602_i2,
  G607_i2,
  G612_i2,
  G617_i2,
  G622_i2,
  G627_i2,
  G632_i2,
  G637_i2,
  n627_lo_buf_i2,
  n639_lo_buf_i2,
  n651_lo_buf_i2,
  n663_lo_buf_i2,
  n675_lo_buf_i2,
  n687_lo_buf_i2,
  n699_lo_buf_i2,
  n711_lo_buf_i2,
  n723_lo_buf_i2,
  n735_lo_buf_i2,
  n747_lo_buf_i2,
  n759_lo_buf_i2,
  n771_lo_buf_i2,
  n783_lo_buf_i2,
  n795_lo_buf_i2,
  n807_lo_buf_i2,
  n819_lo_buf_i2,
  n831_lo_buf_i2,
  n843_lo_buf_i2,
  n855_lo_buf_i2,
  n867_lo_buf_i2,
  n879_lo_buf_i2,
  n891_lo_buf_i2,
  n903_lo_buf_i2,
  n915_lo_buf_i2,
  n927_lo_buf_i2,
  n939_lo_buf_i2,
  n951_lo_buf_i2,
  n963_lo_buf_i2,
  n975_lo_buf_i2,
  n987_lo_buf_i2,
  n999_lo_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input n630_lo;input n642_lo;input n654_lo;input n666_lo;input n678_lo;input n690_lo;input n702_lo;input n714_lo;input n726_lo;input n738_lo;input n750_lo;input n762_lo;input n774_lo;input n786_lo;input n798_lo;input n810_lo;input n822_lo;input n834_lo;input n846_lo;input n858_lo;input n870_lo;input n882_lo;input n894_lo;input n906_lo;input n918_lo;input n930_lo;input n942_lo;input n954_lo;input n966_lo;input n978_lo;input n990_lo;input n1002_lo;input n1005_lo;input n1008_lo;input n1017_lo;input n1020_lo;input n1029_lo;input n1032_lo;input n1041_lo;input n1044_lo;input n1053_lo;input n1056_lo;input n1065_lo;input n1068_lo;input n1077_lo;input n1080_lo;input n1089_lo;input n1092_lo;input n1101_lo;input n1104_lo;input n1837_o2;input n1838_o2;input n1839_o2;input n1840_o2;input n1841_o2;input n1842_o2;input n1843_o2;input n1844_o2;input n1845_o2;input n1846_o2;input n1847_o2;input n1848_o2;input n1849_o2;input n1850_o2;input n1851_o2;input n1852_o2;input n1853_o2;input n1854_o2;input n1855_o2;input n1856_o2;input n1857_o2;input n1858_o2;input n1859_o2;input n1860_o2;input n1861_o2;input n1862_o2;input n1863_o2;input n1864_o2;input n1865_o2;input n1866_o2;input n1867_o2;input n1868_o2;input G834_o2;input G847_o2;input G860_o2;input G873_o2;input G925_o2;input G886_o2;input G912_o2;input G899_o2;input n2151_o2;input n2152_o2;input n2153_o2;input n2154_o2;input n2155_o2;input n2156_o2;input n2157_o2;input n2158_o2;input n2159_o2;input n2160_o2;input n2161_o2;input n2162_o2;input n2163_o2;input n2164_o2;input n2165_o2;input n2166_o2;input n2167_o2;input n2168_o2;input n2169_o2;input n2170_o2;input n2171_o2;input n2172_o2;input n2173_o2;input n2174_o2;input n2175_o2;input n2176_o2;input n2177_o2;input n2178_o2;input n2179_o2;input n2180_o2;input n2181_o2;input n2182_o2;input G974_o2;input G976_o2;input G970_o2;input G972_o2;input G973_o2;input G977_o2;input G971_o2;input G975_o2;input G954_o2;input G956_o2;input G950_o2;input G952_o2;input G953_o2;input G957_o2;input G951_o2;input G955_o2;input G986_o2;input G991_o2;input G770_o2;input G773_o2;input G776_o2;input G779_o2;input G782_o2;input G785_o2;input G788_o2;input G791_o2;input G642_o2;input G645_o2;input G648_o2;input G651_o2;input G654_o2;input G657_o2;input G660_o2;input G663_o2;input G602_o2;input G607_o2;input G612_o2;input G617_o2;input G622_o2;input G627_o2;input G632_o2;input G637_o2;input n627_lo_buf_o2;input n639_lo_buf_o2;input n651_lo_buf_o2;input n663_lo_buf_o2;input n675_lo_buf_o2;input n687_lo_buf_o2;input n699_lo_buf_o2;input n711_lo_buf_o2;input n723_lo_buf_o2;input n735_lo_buf_o2;input n747_lo_buf_o2;input n759_lo_buf_o2;input n771_lo_buf_o2;input n783_lo_buf_o2;input n795_lo_buf_o2;input n807_lo_buf_o2;input n819_lo_buf_o2;input n831_lo_buf_o2;input n843_lo_buf_o2;input n855_lo_buf_o2;input n867_lo_buf_o2;input n879_lo_buf_o2;input n891_lo_buf_o2;input n903_lo_buf_o2;input n915_lo_buf_o2;input n927_lo_buf_o2;input n939_lo_buf_o2;input n951_lo_buf_o2;input n963_lo_buf_o2;input n975_lo_buf_o2;input n987_lo_buf_o2;input n999_lo_buf_o2;
  output G1324;output G1325;output G1326;output G1327;output G1328;output G1329;output G1330;output G1331;output G1332;output G1333;output G1334;output G1335;output G1336;output G1337;output G1338;output G1339;output G1340;output G1341;output G1342;output G1343;output G1344;output G1345;output G1346;output G1347;output G1348;output G1349;output G1350;output G1351;output G1352;output G1353;output G1354;output G1355;output n630_li;output n642_li;output n654_li;output n666_li;output n678_li;output n690_li;output n702_li;output n714_li;output n726_li;output n738_li;output n750_li;output n762_li;output n774_li;output n786_li;output n798_li;output n810_li;output n822_li;output n834_li;output n846_li;output n858_li;output n870_li;output n882_li;output n894_li;output n906_li;output n918_li;output n930_li;output n942_li;output n954_li;output n966_li;output n978_li;output n990_li;output n1002_li;output n1005_li;output n1008_li;output n1017_li;output n1020_li;output n1029_li;output n1032_li;output n1041_li;output n1044_li;output n1053_li;output n1056_li;output n1065_li;output n1068_li;output n1077_li;output n1080_li;output n1089_li;output n1092_li;output n1101_li;output n1104_li;output n1837_i2;output n1838_i2;output n1839_i2;output n1840_i2;output n1841_i2;output n1842_i2;output n1843_i2;output n1844_i2;output n1845_i2;output n1846_i2;output n1847_i2;output n1848_i2;output n1849_i2;output n1850_i2;output n1851_i2;output n1852_i2;output n1853_i2;output n1854_i2;output n1855_i2;output n1856_i2;output n1857_i2;output n1858_i2;output n1859_i2;output n1860_i2;output n1861_i2;output n1862_i2;output n1863_i2;output n1864_i2;output n1865_i2;output n1866_i2;output n1867_i2;output n1868_i2;output G834_i2;output G847_i2;output G860_i2;output G873_i2;output G925_i2;output G886_i2;output G912_i2;output G899_i2;output n2151_i2;output n2152_i2;output n2153_i2;output n2154_i2;output n2155_i2;output n2156_i2;output n2157_i2;output n2158_i2;output n2159_i2;output n2160_i2;output n2161_i2;output n2162_i2;output n2163_i2;output n2164_i2;output n2165_i2;output n2166_i2;output n2167_i2;output n2168_i2;output n2169_i2;output n2170_i2;output n2171_i2;output n2172_i2;output n2173_i2;output n2174_i2;output n2175_i2;output n2176_i2;output n2177_i2;output n2178_i2;output n2179_i2;output n2180_i2;output n2181_i2;output n2182_i2;output G974_i2;output G976_i2;output G970_i2;output G972_i2;output G973_i2;output G977_i2;output G971_i2;output G975_i2;output G954_i2;output G956_i2;output G950_i2;output G952_i2;output G953_i2;output G957_i2;output G951_i2;output G955_i2;output G986_i2;output G991_i2;output G770_i2;output G773_i2;output G776_i2;output G779_i2;output G782_i2;output G785_i2;output G788_i2;output G791_i2;output G642_i2;output G645_i2;output G648_i2;output G651_i2;output G654_i2;output G657_i2;output G660_i2;output G663_i2;output G602_i2;output G607_i2;output G612_i2;output G617_i2;output G622_i2;output G627_i2;output G632_i2;output G637_i2;output n627_lo_buf_i2;output n639_lo_buf_i2;output n651_lo_buf_i2;output n663_lo_buf_i2;output n675_lo_buf_i2;output n687_lo_buf_i2;output n699_lo_buf_i2;output n711_lo_buf_i2;output n723_lo_buf_i2;output n735_lo_buf_i2;output n747_lo_buf_i2;output n759_lo_buf_i2;output n771_lo_buf_i2;output n783_lo_buf_i2;output n795_lo_buf_i2;output n807_lo_buf_i2;output n819_lo_buf_i2;output n831_lo_buf_i2;output n843_lo_buf_i2;output n855_lo_buf_i2;output n867_lo_buf_i2;output n879_lo_buf_i2;output n891_lo_buf_i2;output n903_lo_buf_i2;output n915_lo_buf_i2;output n927_lo_buf_i2;output n939_lo_buf_i2;output n951_lo_buf_i2;output n963_lo_buf_i2;output n975_lo_buf_i2;output n987_lo_buf_i2;output n999_lo_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire n630_lo_p;
  wire n630_lo_n;
  wire n642_lo_p;
  wire n642_lo_n;
  wire n654_lo_p;
  wire n654_lo_n;
  wire n666_lo_p;
  wire n666_lo_n;
  wire n678_lo_p;
  wire n678_lo_n;
  wire n690_lo_p;
  wire n690_lo_n;
  wire n702_lo_p;
  wire n702_lo_n;
  wire n714_lo_p;
  wire n714_lo_n;
  wire n726_lo_p;
  wire n726_lo_n;
  wire n738_lo_p;
  wire n738_lo_n;
  wire n750_lo_p;
  wire n750_lo_n;
  wire n762_lo_p;
  wire n762_lo_n;
  wire n774_lo_p;
  wire n774_lo_n;
  wire n786_lo_p;
  wire n786_lo_n;
  wire n798_lo_p;
  wire n798_lo_n;
  wire n810_lo_p;
  wire n810_lo_n;
  wire n822_lo_p;
  wire n822_lo_n;
  wire n834_lo_p;
  wire n834_lo_n;
  wire n846_lo_p;
  wire n846_lo_n;
  wire n858_lo_p;
  wire n858_lo_n;
  wire n870_lo_p;
  wire n870_lo_n;
  wire n882_lo_p;
  wire n882_lo_n;
  wire n894_lo_p;
  wire n894_lo_n;
  wire n906_lo_p;
  wire n906_lo_n;
  wire n918_lo_p;
  wire n918_lo_n;
  wire n930_lo_p;
  wire n930_lo_n;
  wire n942_lo_p;
  wire n942_lo_n;
  wire n954_lo_p;
  wire n954_lo_n;
  wire n966_lo_p;
  wire n966_lo_n;
  wire n978_lo_p;
  wire n978_lo_n;
  wire n990_lo_p;
  wire n990_lo_n;
  wire n1002_lo_p;
  wire n1002_lo_n;
  wire n1005_lo_p;
  wire n1005_lo_n;
  wire n1008_lo_p;
  wire n1008_lo_n;
  wire n1017_lo_p;
  wire n1017_lo_n;
  wire n1020_lo_p;
  wire n1020_lo_n;
  wire n1029_lo_p;
  wire n1029_lo_n;
  wire n1032_lo_p;
  wire n1032_lo_n;
  wire n1041_lo_p;
  wire n1041_lo_n;
  wire n1044_lo_p;
  wire n1044_lo_n;
  wire n1053_lo_p;
  wire n1053_lo_n;
  wire n1056_lo_p;
  wire n1056_lo_n;
  wire n1065_lo_p;
  wire n1065_lo_n;
  wire n1068_lo_p;
  wire n1068_lo_n;
  wire n1077_lo_p;
  wire n1077_lo_n;
  wire n1080_lo_p;
  wire n1080_lo_n;
  wire n1089_lo_p;
  wire n1089_lo_n;
  wire n1092_lo_p;
  wire n1092_lo_n;
  wire n1101_lo_p;
  wire n1101_lo_n;
  wire n1104_lo_p;
  wire n1104_lo_n;
  wire n1837_o2_p;
  wire n1837_o2_n;
  wire n1838_o2_p;
  wire n1838_o2_n;
  wire n1839_o2_p;
  wire n1839_o2_n;
  wire n1840_o2_p;
  wire n1840_o2_n;
  wire n1841_o2_p;
  wire n1841_o2_n;
  wire n1842_o2_p;
  wire n1842_o2_n;
  wire n1843_o2_p;
  wire n1843_o2_n;
  wire n1844_o2_p;
  wire n1844_o2_n;
  wire n1845_o2_p;
  wire n1845_o2_n;
  wire n1846_o2_p;
  wire n1846_o2_n;
  wire n1847_o2_p;
  wire n1847_o2_n;
  wire n1848_o2_p;
  wire n1848_o2_n;
  wire n1849_o2_p;
  wire n1849_o2_n;
  wire n1850_o2_p;
  wire n1850_o2_n;
  wire n1851_o2_p;
  wire n1851_o2_n;
  wire n1852_o2_p;
  wire n1852_o2_n;
  wire n1853_o2_p;
  wire n1853_o2_n;
  wire n1854_o2_p;
  wire n1854_o2_n;
  wire n1855_o2_p;
  wire n1855_o2_n;
  wire n1856_o2_p;
  wire n1856_o2_n;
  wire n1857_o2_p;
  wire n1857_o2_n;
  wire n1858_o2_p;
  wire n1858_o2_n;
  wire n1859_o2_p;
  wire n1859_o2_n;
  wire n1860_o2_p;
  wire n1860_o2_n;
  wire n1861_o2_p;
  wire n1861_o2_n;
  wire n1862_o2_p;
  wire n1862_o2_n;
  wire n1863_o2_p;
  wire n1863_o2_n;
  wire n1864_o2_p;
  wire n1864_o2_n;
  wire n1865_o2_p;
  wire n1865_o2_n;
  wire n1866_o2_p;
  wire n1866_o2_n;
  wire n1867_o2_p;
  wire n1867_o2_n;
  wire n1868_o2_p;
  wire n1868_o2_n;
  wire G834_o2_p;
  wire G834_o2_n;
  wire G847_o2_p;
  wire G847_o2_n;
  wire G860_o2_p;
  wire G860_o2_n;
  wire G873_o2_p;
  wire G873_o2_n;
  wire G925_o2_p;
  wire G925_o2_n;
  wire G886_o2_p;
  wire G886_o2_n;
  wire G912_o2_p;
  wire G912_o2_n;
  wire G899_o2_p;
  wire G899_o2_n;
  wire n2151_o2_p;
  wire n2151_o2_n;
  wire n2152_o2_p;
  wire n2152_o2_n;
  wire n2153_o2_p;
  wire n2153_o2_n;
  wire n2154_o2_p;
  wire n2154_o2_n;
  wire n2155_o2_p;
  wire n2155_o2_n;
  wire n2156_o2_p;
  wire n2156_o2_n;
  wire n2157_o2_p;
  wire n2157_o2_n;
  wire n2158_o2_p;
  wire n2158_o2_n;
  wire n2159_o2_p;
  wire n2159_o2_n;
  wire n2160_o2_p;
  wire n2160_o2_n;
  wire n2161_o2_p;
  wire n2161_o2_n;
  wire n2162_o2_p;
  wire n2162_o2_n;
  wire n2163_o2_p;
  wire n2163_o2_n;
  wire n2164_o2_p;
  wire n2164_o2_n;
  wire n2165_o2_p;
  wire n2165_o2_n;
  wire n2166_o2_p;
  wire n2166_o2_n;
  wire n2167_o2_p;
  wire n2167_o2_n;
  wire n2168_o2_p;
  wire n2168_o2_n;
  wire n2169_o2_p;
  wire n2169_o2_n;
  wire n2170_o2_p;
  wire n2170_o2_n;
  wire n2171_o2_p;
  wire n2171_o2_n;
  wire n2172_o2_p;
  wire n2172_o2_n;
  wire n2173_o2_p;
  wire n2173_o2_n;
  wire n2174_o2_p;
  wire n2174_o2_n;
  wire n2175_o2_p;
  wire n2175_o2_n;
  wire n2176_o2_p;
  wire n2176_o2_n;
  wire n2177_o2_p;
  wire n2177_o2_n;
  wire n2178_o2_p;
  wire n2178_o2_n;
  wire n2179_o2_p;
  wire n2179_o2_n;
  wire n2180_o2_p;
  wire n2180_o2_n;
  wire n2181_o2_p;
  wire n2181_o2_n;
  wire n2182_o2_p;
  wire n2182_o2_n;
  wire G974_o2_p;
  wire G974_o2_n;
  wire G976_o2_p;
  wire G976_o2_n;
  wire G970_o2_p;
  wire G970_o2_n;
  wire G972_o2_p;
  wire G972_o2_n;
  wire G973_o2_p;
  wire G973_o2_n;
  wire G977_o2_p;
  wire G977_o2_n;
  wire G971_o2_p;
  wire G971_o2_n;
  wire G975_o2_p;
  wire G975_o2_n;
  wire G954_o2_p;
  wire G954_o2_n;
  wire G956_o2_p;
  wire G956_o2_n;
  wire G950_o2_p;
  wire G950_o2_n;
  wire G952_o2_p;
  wire G952_o2_n;
  wire G953_o2_p;
  wire G953_o2_n;
  wire G957_o2_p;
  wire G957_o2_n;
  wire G951_o2_p;
  wire G951_o2_n;
  wire G955_o2_p;
  wire G955_o2_n;
  wire G986_o2_p;
  wire G986_o2_n;
  wire G991_o2_p;
  wire G991_o2_n;
  wire G770_o2_p;
  wire G770_o2_n;
  wire G773_o2_p;
  wire G773_o2_n;
  wire G776_o2_p;
  wire G776_o2_n;
  wire G779_o2_p;
  wire G779_o2_n;
  wire G782_o2_p;
  wire G782_o2_n;
  wire G785_o2_p;
  wire G785_o2_n;
  wire G788_o2_p;
  wire G788_o2_n;
  wire G791_o2_p;
  wire G791_o2_n;
  wire G642_o2_p;
  wire G642_o2_n;
  wire G645_o2_p;
  wire G645_o2_n;
  wire G648_o2_p;
  wire G648_o2_n;
  wire G651_o2_p;
  wire G651_o2_n;
  wire G654_o2_p;
  wire G654_o2_n;
  wire G657_o2_p;
  wire G657_o2_n;
  wire G660_o2_p;
  wire G660_o2_n;
  wire G663_o2_p;
  wire G663_o2_n;
  wire G602_o2_p;
  wire G602_o2_n;
  wire G607_o2_p;
  wire G607_o2_n;
  wire G612_o2_p;
  wire G612_o2_n;
  wire G617_o2_p;
  wire G617_o2_n;
  wire G622_o2_p;
  wire G622_o2_n;
  wire G627_o2_p;
  wire G627_o2_n;
  wire G632_o2_p;
  wire G632_o2_n;
  wire G637_o2_p;
  wire G637_o2_n;
  wire n627_lo_buf_o2_p;
  wire n627_lo_buf_o2_n;
  wire n639_lo_buf_o2_p;
  wire n639_lo_buf_o2_n;
  wire n651_lo_buf_o2_p;
  wire n651_lo_buf_o2_n;
  wire n663_lo_buf_o2_p;
  wire n663_lo_buf_o2_n;
  wire n675_lo_buf_o2_p;
  wire n675_lo_buf_o2_n;
  wire n687_lo_buf_o2_p;
  wire n687_lo_buf_o2_n;
  wire n699_lo_buf_o2_p;
  wire n699_lo_buf_o2_n;
  wire n711_lo_buf_o2_p;
  wire n711_lo_buf_o2_n;
  wire n723_lo_buf_o2_p;
  wire n723_lo_buf_o2_n;
  wire n735_lo_buf_o2_p;
  wire n735_lo_buf_o2_n;
  wire n747_lo_buf_o2_p;
  wire n747_lo_buf_o2_n;
  wire n759_lo_buf_o2_p;
  wire n759_lo_buf_o2_n;
  wire n771_lo_buf_o2_p;
  wire n771_lo_buf_o2_n;
  wire n783_lo_buf_o2_p;
  wire n783_lo_buf_o2_n;
  wire n795_lo_buf_o2_p;
  wire n795_lo_buf_o2_n;
  wire n807_lo_buf_o2_p;
  wire n807_lo_buf_o2_n;
  wire n819_lo_buf_o2_p;
  wire n819_lo_buf_o2_n;
  wire n831_lo_buf_o2_p;
  wire n831_lo_buf_o2_n;
  wire n843_lo_buf_o2_p;
  wire n843_lo_buf_o2_n;
  wire n855_lo_buf_o2_p;
  wire n855_lo_buf_o2_n;
  wire n867_lo_buf_o2_p;
  wire n867_lo_buf_o2_n;
  wire n879_lo_buf_o2_p;
  wire n879_lo_buf_o2_n;
  wire n891_lo_buf_o2_p;
  wire n891_lo_buf_o2_n;
  wire n903_lo_buf_o2_p;
  wire n903_lo_buf_o2_n;
  wire n915_lo_buf_o2_p;
  wire n915_lo_buf_o2_n;
  wire n927_lo_buf_o2_p;
  wire n927_lo_buf_o2_n;
  wire n939_lo_buf_o2_p;
  wire n939_lo_buf_o2_n;
  wire n951_lo_buf_o2_p;
  wire n951_lo_buf_o2_n;
  wire n963_lo_buf_o2_p;
  wire n963_lo_buf_o2_n;
  wire n975_lo_buf_o2_p;
  wire n975_lo_buf_o2_n;
  wire n987_lo_buf_o2_p;
  wire n987_lo_buf_o2_n;
  wire n999_lo_buf_o2_p;
  wire n999_lo_buf_o2_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire G925_o2_p_spl_;
  wire G925_o2_p_spl_0;
  wire G925_o2_p_spl_00;
  wire G925_o2_p_spl_01;
  wire G925_o2_p_spl_1;
  wire G925_o2_n_spl_;
  wire G925_o2_n_spl_0;
  wire G925_o2_n_spl_00;
  wire G925_o2_n_spl_01;
  wire G925_o2_n_spl_1;
  wire G912_o2_p_spl_;
  wire G912_o2_p_spl_0;
  wire G912_o2_p_spl_00;
  wire G912_o2_p_spl_01;
  wire G912_o2_p_spl_1;
  wire G912_o2_n_spl_;
  wire G912_o2_n_spl_0;
  wire G912_o2_n_spl_00;
  wire G912_o2_n_spl_01;
  wire G912_o2_n_spl_1;
  wire G986_o2_p_spl_;
  wire G986_o2_p_spl_0;
  wire G986_o2_p_spl_1;
  wire G986_o2_n_spl_;
  wire G986_o2_n_spl_0;
  wire G986_o2_n_spl_1;
  wire g241_p_spl_;
  wire g241_p_spl_0;
  wire g241_p_spl_1;
  wire G834_o2_p_spl_;
  wire G834_o2_p_spl_0;
  wire G834_o2_p_spl_00;
  wire G834_o2_p_spl_01;
  wire G834_o2_p_spl_1;
  wire g241_n_spl_;
  wire g241_n_spl_0;
  wire g241_n_spl_1;
  wire G834_o2_n_spl_;
  wire G834_o2_n_spl_0;
  wire G834_o2_n_spl_00;
  wire G834_o2_n_spl_01;
  wire G834_o2_n_spl_1;
  wire g243_n_spl_;
  wire G847_o2_p_spl_;
  wire G847_o2_p_spl_0;
  wire G847_o2_p_spl_00;
  wire G847_o2_p_spl_01;
  wire G847_o2_p_spl_1;
  wire G847_o2_n_spl_;
  wire G847_o2_n_spl_0;
  wire G847_o2_n_spl_00;
  wire G847_o2_n_spl_01;
  wire G847_o2_n_spl_1;
  wire g248_n_spl_;
  wire G860_o2_p_spl_;
  wire G860_o2_p_spl_0;
  wire G860_o2_p_spl_00;
  wire G860_o2_p_spl_01;
  wire G860_o2_p_spl_1;
  wire G860_o2_n_spl_;
  wire G860_o2_n_spl_0;
  wire G860_o2_n_spl_00;
  wire G860_o2_n_spl_01;
  wire G860_o2_n_spl_1;
  wire g253_n_spl_;
  wire G873_o2_p_spl_;
  wire G873_o2_p_spl_0;
  wire G873_o2_p_spl_00;
  wire G873_o2_p_spl_01;
  wire G873_o2_p_spl_1;
  wire G873_o2_n_spl_;
  wire G873_o2_n_spl_0;
  wire G873_o2_n_spl_00;
  wire G873_o2_n_spl_01;
  wire G873_o2_n_spl_1;
  wire g258_n_spl_;
  wire G899_o2_p_spl_;
  wire G899_o2_p_spl_0;
  wire G899_o2_p_spl_00;
  wire G899_o2_p_spl_01;
  wire G899_o2_p_spl_1;
  wire G899_o2_n_spl_;
  wire G899_o2_n_spl_0;
  wire G899_o2_n_spl_00;
  wire G899_o2_n_spl_01;
  wire G899_o2_n_spl_1;
  wire g265_p_spl_;
  wire g265_p_spl_0;
  wire g265_p_spl_1;
  wire g265_n_spl_;
  wire g265_n_spl_0;
  wire g265_n_spl_1;
  wire g267_n_spl_;
  wire g272_n_spl_;
  wire g277_n_spl_;
  wire g282_n_spl_;
  wire G886_o2_p_spl_;
  wire G886_o2_p_spl_0;
  wire G886_o2_p_spl_00;
  wire G886_o2_p_spl_01;
  wire G886_o2_p_spl_1;
  wire G886_o2_n_spl_;
  wire G886_o2_n_spl_0;
  wire G886_o2_n_spl_00;
  wire G886_o2_n_spl_01;
  wire G886_o2_n_spl_1;
  wire g289_p_spl_;
  wire g289_p_spl_0;
  wire g289_p_spl_1;
  wire g289_n_spl_;
  wire g289_n_spl_0;
  wire g289_n_spl_1;
  wire g291_n_spl_;
  wire g296_n_spl_;
  wire g301_n_spl_;
  wire g306_n_spl_;
  wire g313_p_spl_;
  wire g313_p_spl_0;
  wire g313_p_spl_1;
  wire g313_n_spl_;
  wire g313_n_spl_0;
  wire g313_n_spl_1;
  wire g315_n_spl_;
  wire g320_n_spl_;
  wire g325_n_spl_;
  wire g330_n_spl_;
  wire G991_o2_p_spl_;
  wire G991_o2_p_spl_0;
  wire G991_o2_p_spl_1;
  wire G991_o2_n_spl_;
  wire G991_o2_n_spl_0;
  wire G991_o2_n_spl_1;
  wire g337_p_spl_;
  wire g337_p_spl_0;
  wire g337_p_spl_1;
  wire g337_n_spl_;
  wire g337_n_spl_0;
  wire g337_n_spl_1;
  wire g339_n_spl_;
  wire g344_n_spl_;
  wire g349_n_spl_;
  wire g354_n_spl_;
  wire g361_p_spl_;
  wire g361_p_spl_0;
  wire g361_p_spl_1;
  wire g361_n_spl_;
  wire g361_n_spl_0;
  wire g361_n_spl_1;
  wire g363_n_spl_;
  wire g368_n_spl_;
  wire g373_n_spl_;
  wire g378_n_spl_;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g385_p_spl_1;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g385_n_spl_1;
  wire g387_n_spl_;
  wire g392_n_spl_;
  wire g397_n_spl_;
  wire g402_n_spl_;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g409_p_spl_1;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g409_n_spl_1;
  wire g411_n_spl_;
  wire g416_n_spl_;
  wire g421_n_spl_;
  wire g426_n_spl_;
  wire G642_o2_p_spl_;
  wire G770_o2_p_spl_;
  wire G642_o2_n_spl_;
  wire G770_o2_n_spl_;
  wire g430_n_spl_;
  wire g430_p_spl_;
  wire G645_o2_p_spl_;
  wire G773_o2_p_spl_;
  wire G645_o2_n_spl_;
  wire G773_o2_n_spl_;
  wire g434_n_spl_;
  wire g434_p_spl_;
  wire G648_o2_p_spl_;
  wire G776_o2_p_spl_;
  wire G648_o2_n_spl_;
  wire G776_o2_n_spl_;
  wire g438_n_spl_;
  wire g438_p_spl_;
  wire G651_o2_p_spl_;
  wire G779_o2_p_spl_;
  wire G651_o2_n_spl_;
  wire G779_o2_n_spl_;
  wire g442_n_spl_;
  wire g442_p_spl_;
  wire G654_o2_p_spl_;
  wire G782_o2_p_spl_;
  wire G654_o2_n_spl_;
  wire G782_o2_n_spl_;
  wire g446_n_spl_;
  wire g446_p_spl_;
  wire G657_o2_p_spl_;
  wire G785_o2_p_spl_;
  wire G657_o2_n_spl_;
  wire G785_o2_n_spl_;
  wire g450_n_spl_;
  wire g450_p_spl_;
  wire G660_o2_p_spl_;
  wire G788_o2_p_spl_;
  wire G660_o2_n_spl_;
  wire G788_o2_n_spl_;
  wire g454_n_spl_;
  wire g454_p_spl_;
  wire G663_o2_p_spl_;
  wire G791_o2_p_spl_;
  wire G663_o2_n_spl_;
  wire G791_o2_n_spl_;
  wire g458_n_spl_;
  wire g458_p_spl_;
  wire g437_n_spl_;
  wire g433_n_spl_;
  wire g462_n_spl_;
  wire g441_n_spl_;
  wire g441_n_spl_0;
  wire g445_p_spl_;
  wire g445_p_spl_0;
  wire g445_p_spl_1;
  wire g441_p_spl_;
  wire g441_p_spl_0;
  wire g441_p_spl_1;
  wire g445_n_spl_;
  wire g445_n_spl_0;
  wire g437_p_spl_;
  wire g437_p_spl_0;
  wire g437_p_spl_1;
  wire g433_p_spl_;
  wire g433_p_spl_0;
  wire g433_p_spl_1;
  wire g453_n_spl_;
  wire g449_n_spl_;
  wire g476_n_spl_;
  wire g457_n_spl_;
  wire g457_n_spl_0;
  wire g461_p_spl_;
  wire g461_p_spl_0;
  wire g461_p_spl_1;
  wire g457_p_spl_;
  wire g457_p_spl_0;
  wire g457_p_spl_1;
  wire g461_n_spl_;
  wire g461_n_spl_0;
  wire g453_p_spl_;
  wire g453_p_spl_0;
  wire g453_p_spl_1;
  wire g449_p_spl_;
  wire g449_p_spl_0;
  wire g449_p_spl_1;
  wire n1104_lo_p_spl_;
  wire n1104_lo_p_spl_0;
  wire n1104_lo_p_spl_00;
  wire n1104_lo_p_spl_01;
  wire n1104_lo_p_spl_1;
  wire n1104_lo_p_spl_10;
  wire n1104_lo_p_spl_11;
  wire n1104_lo_n_spl_;
  wire n1104_lo_n_spl_0;
  wire n1104_lo_n_spl_00;
  wire n1104_lo_n_spl_01;
  wire n1104_lo_n_spl_1;
  wire n1104_lo_n_spl_10;
  wire n1104_lo_n_spl_11;
  wire G627_o2_p_spl_;
  wire G627_o2_p_spl_0;
  wire G627_o2_p_spl_1;
  wire G622_o2_p_spl_;
  wire G622_o2_p_spl_0;
  wire G622_o2_p_spl_1;
  wire G627_o2_n_spl_;
  wire G627_o2_n_spl_0;
  wire G627_o2_n_spl_1;
  wire G622_o2_n_spl_;
  wire G622_o2_n_spl_0;
  wire G622_o2_n_spl_1;
  wire g491_n_spl_;
  wire g491_p_spl_;
  wire g495_p_spl_;
  wire G637_o2_p_spl_;
  wire G637_o2_p_spl_0;
  wire G637_o2_p_spl_1;
  wire G632_o2_p_spl_;
  wire G632_o2_p_spl_0;
  wire G632_o2_p_spl_1;
  wire G637_o2_n_spl_;
  wire G637_o2_n_spl_0;
  wire G637_o2_n_spl_1;
  wire G632_o2_n_spl_;
  wire G632_o2_n_spl_0;
  wire G632_o2_n_spl_1;
  wire g500_n_spl_;
  wire g500_p_spl_;
  wire g504_p_spl_;
  wire g509_n_spl_;
  wire g509_p_spl_;
  wire g513_p_spl_;
  wire g518_n_spl_;
  wire g518_p_spl_;
  wire g522_p_spl_;
  wire G607_o2_p_spl_;
  wire G607_o2_p_spl_0;
  wire G607_o2_p_spl_1;
  wire G602_o2_p_spl_;
  wire G602_o2_p_spl_0;
  wire G602_o2_p_spl_1;
  wire G607_o2_n_spl_;
  wire G607_o2_n_spl_0;
  wire G607_o2_n_spl_1;
  wire G602_o2_n_spl_;
  wire G602_o2_n_spl_0;
  wire G602_o2_n_spl_1;
  wire g527_n_spl_;
  wire g527_p_spl_;
  wire g531_p_spl_;
  wire G617_o2_p_spl_;
  wire G617_o2_p_spl_0;
  wire G617_o2_p_spl_1;
  wire G612_o2_p_spl_;
  wire G612_o2_p_spl_0;
  wire G612_o2_p_spl_1;
  wire G617_o2_n_spl_;
  wire G617_o2_n_spl_0;
  wire G617_o2_n_spl_1;
  wire G612_o2_n_spl_;
  wire G612_o2_n_spl_0;
  wire G612_o2_n_spl_1;
  wire g536_n_spl_;
  wire g536_p_spl_;
  wire g540_p_spl_;
  wire g545_n_spl_;
  wire g545_p_spl_;
  wire g549_p_spl_;
  wire g554_n_spl_;
  wire g554_p_spl_;
  wire g558_p_spl_;
  wire n2155_o2_p_spl_;
  wire n2151_o2_p_spl_;
  wire n2155_o2_n_spl_;
  wire n2155_o2_n_spl_0;
  wire n2151_o2_n_spl_;
  wire n2151_o2_n_spl_0;
  wire g562_n_spl_;
  wire g562_p_spl_;
  wire n2163_o2_p_spl_;
  wire n2159_o2_p_spl_;
  wire n2163_o2_n_spl_;
  wire n2163_o2_n_spl_0;
  wire n2159_o2_n_spl_;
  wire n2159_o2_n_spl_0;
  wire g566_n_spl_;
  wire g566_p_spl_;
  wire g570_p_spl_;
  wire n2156_o2_p_spl_;
  wire n2152_o2_p_spl_;
  wire n2156_o2_n_spl_;
  wire n2156_o2_n_spl_0;
  wire n2152_o2_n_spl_;
  wire n2152_o2_n_spl_0;
  wire g574_n_spl_;
  wire g574_p_spl_;
  wire n2164_o2_p_spl_;
  wire n2160_o2_p_spl_;
  wire n2164_o2_n_spl_;
  wire n2164_o2_n_spl_0;
  wire n2160_o2_n_spl_;
  wire n2160_o2_n_spl_0;
  wire g578_n_spl_;
  wire g578_p_spl_;
  wire g582_p_spl_;
  wire n2157_o2_p_spl_;
  wire n2153_o2_p_spl_;
  wire n2157_o2_n_spl_;
  wire n2157_o2_n_spl_0;
  wire n2153_o2_n_spl_;
  wire n2153_o2_n_spl_0;
  wire g586_n_spl_;
  wire g586_p_spl_;
  wire n2165_o2_p_spl_;
  wire n2161_o2_p_spl_;
  wire n2165_o2_n_spl_;
  wire n2165_o2_n_spl_0;
  wire n2161_o2_n_spl_;
  wire n2161_o2_n_spl_0;
  wire g590_n_spl_;
  wire g590_p_spl_;
  wire g594_p_spl_;
  wire n2158_o2_p_spl_;
  wire n2154_o2_p_spl_;
  wire n2158_o2_n_spl_;
  wire n2158_o2_n_spl_0;
  wire n2154_o2_n_spl_;
  wire n2154_o2_n_spl_0;
  wire g598_n_spl_;
  wire g598_p_spl_;
  wire n2166_o2_p_spl_;
  wire n2162_o2_p_spl_;
  wire n2166_o2_n_spl_;
  wire n2166_o2_n_spl_0;
  wire n2162_o2_n_spl_;
  wire n2162_o2_n_spl_0;
  wire g602_n_spl_;
  wire g602_p_spl_;
  wire g606_p_spl_;
  wire n2171_o2_p_spl_;
  wire n2167_o2_p_spl_;
  wire n2171_o2_n_spl_;
  wire n2171_o2_n_spl_0;
  wire n2167_o2_n_spl_;
  wire n2167_o2_n_spl_0;
  wire g610_n_spl_;
  wire g610_p_spl_;
  wire n2179_o2_p_spl_;
  wire n2175_o2_p_spl_;
  wire n2179_o2_n_spl_;
  wire n2179_o2_n_spl_0;
  wire n2175_o2_n_spl_;
  wire n2175_o2_n_spl_0;
  wire g614_n_spl_;
  wire g614_p_spl_;
  wire g618_p_spl_;
  wire n2172_o2_p_spl_;
  wire n2168_o2_p_spl_;
  wire n2172_o2_n_spl_;
  wire n2172_o2_n_spl_0;
  wire n2168_o2_n_spl_;
  wire n2168_o2_n_spl_0;
  wire g622_n_spl_;
  wire g622_p_spl_;
  wire n2180_o2_p_spl_;
  wire n2176_o2_p_spl_;
  wire n2180_o2_n_spl_;
  wire n2180_o2_n_spl_0;
  wire n2176_o2_n_spl_;
  wire n2176_o2_n_spl_0;
  wire g626_n_spl_;
  wire g626_p_spl_;
  wire g630_p_spl_;
  wire n2173_o2_p_spl_;
  wire n2169_o2_p_spl_;
  wire n2173_o2_n_spl_;
  wire n2173_o2_n_spl_0;
  wire n2169_o2_n_spl_;
  wire n2169_o2_n_spl_0;
  wire g634_n_spl_;
  wire g634_p_spl_;
  wire n2181_o2_p_spl_;
  wire n2177_o2_p_spl_;
  wire n2181_o2_n_spl_;
  wire n2181_o2_n_spl_0;
  wire n2177_o2_n_spl_;
  wire n2177_o2_n_spl_0;
  wire g638_n_spl_;
  wire g638_p_spl_;
  wire g642_p_spl_;
  wire n2174_o2_p_spl_;
  wire n2170_o2_p_spl_;
  wire n2174_o2_n_spl_;
  wire n2174_o2_n_spl_0;
  wire n2170_o2_n_spl_;
  wire n2170_o2_n_spl_0;
  wire g646_n_spl_;
  wire g646_p_spl_;
  wire n2182_o2_p_spl_;
  wire n2178_o2_p_spl_;
  wire n2182_o2_n_spl_;
  wire n2182_o2_n_spl_0;
  wire n2178_o2_n_spl_;
  wire n2178_o2_n_spl_0;
  wire g650_n_spl_;
  wire g650_p_spl_;
  wire g654_p_spl_;
  wire n639_lo_buf_o2_p_spl_;
  wire n627_lo_buf_o2_p_spl_;
  wire n639_lo_buf_o2_n_spl_;
  wire n639_lo_buf_o2_n_spl_0;
  wire n627_lo_buf_o2_n_spl_;
  wire n627_lo_buf_o2_n_spl_0;
  wire g658_n_spl_;
  wire g658_p_spl_;
  wire n663_lo_buf_o2_p_spl_;
  wire n651_lo_buf_o2_p_spl_;
  wire n663_lo_buf_o2_n_spl_;
  wire n663_lo_buf_o2_n_spl_0;
  wire n651_lo_buf_o2_n_spl_;
  wire n651_lo_buf_o2_n_spl_0;
  wire g662_n_spl_;
  wire g662_p_spl_;
  wire g666_p_spl_;
  wire n687_lo_buf_o2_p_spl_;
  wire n675_lo_buf_o2_p_spl_;
  wire n687_lo_buf_o2_n_spl_;
  wire n687_lo_buf_o2_n_spl_0;
  wire n675_lo_buf_o2_n_spl_;
  wire n675_lo_buf_o2_n_spl_0;
  wire g670_n_spl_;
  wire g670_p_spl_;
  wire n711_lo_buf_o2_p_spl_;
  wire n699_lo_buf_o2_p_spl_;
  wire n711_lo_buf_o2_n_spl_;
  wire n711_lo_buf_o2_n_spl_0;
  wire n699_lo_buf_o2_n_spl_;
  wire n699_lo_buf_o2_n_spl_0;
  wire g674_n_spl_;
  wire g674_p_spl_;
  wire g678_p_spl_;
  wire n735_lo_buf_o2_p_spl_;
  wire n723_lo_buf_o2_p_spl_;
  wire n735_lo_buf_o2_n_spl_;
  wire n735_lo_buf_o2_n_spl_0;
  wire n723_lo_buf_o2_n_spl_;
  wire n723_lo_buf_o2_n_spl_0;
  wire g682_n_spl_;
  wire g682_p_spl_;
  wire n759_lo_buf_o2_p_spl_;
  wire n747_lo_buf_o2_p_spl_;
  wire n759_lo_buf_o2_n_spl_;
  wire n759_lo_buf_o2_n_spl_0;
  wire n747_lo_buf_o2_n_spl_;
  wire n747_lo_buf_o2_n_spl_0;
  wire g686_n_spl_;
  wire g686_p_spl_;
  wire g690_p_spl_;
  wire n783_lo_buf_o2_p_spl_;
  wire n771_lo_buf_o2_p_spl_;
  wire n783_lo_buf_o2_n_spl_;
  wire n783_lo_buf_o2_n_spl_0;
  wire n771_lo_buf_o2_n_spl_;
  wire n771_lo_buf_o2_n_spl_0;
  wire g694_n_spl_;
  wire g694_p_spl_;
  wire n807_lo_buf_o2_p_spl_;
  wire n795_lo_buf_o2_p_spl_;
  wire n807_lo_buf_o2_n_spl_;
  wire n807_lo_buf_o2_n_spl_0;
  wire n795_lo_buf_o2_n_spl_;
  wire n795_lo_buf_o2_n_spl_0;
  wire g698_n_spl_;
  wire g698_p_spl_;
  wire g702_p_spl_;
  wire n831_lo_buf_o2_p_spl_;
  wire n819_lo_buf_o2_p_spl_;
  wire n831_lo_buf_o2_n_spl_;
  wire n831_lo_buf_o2_n_spl_0;
  wire n819_lo_buf_o2_n_spl_;
  wire n819_lo_buf_o2_n_spl_0;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire n855_lo_buf_o2_p_spl_;
  wire n843_lo_buf_o2_p_spl_;
  wire n855_lo_buf_o2_n_spl_;
  wire n855_lo_buf_o2_n_spl_0;
  wire n843_lo_buf_o2_n_spl_;
  wire n843_lo_buf_o2_n_spl_0;
  wire g710_n_spl_;
  wire g710_p_spl_;
  wire g714_p_spl_;
  wire n879_lo_buf_o2_p_spl_;
  wire n867_lo_buf_o2_p_spl_;
  wire n879_lo_buf_o2_n_spl_;
  wire n879_lo_buf_o2_n_spl_0;
  wire n867_lo_buf_o2_n_spl_;
  wire n867_lo_buf_o2_n_spl_0;
  wire g718_n_spl_;
  wire g718_p_spl_;
  wire n903_lo_buf_o2_p_spl_;
  wire n891_lo_buf_o2_p_spl_;
  wire n903_lo_buf_o2_n_spl_;
  wire n903_lo_buf_o2_n_spl_0;
  wire n891_lo_buf_o2_n_spl_;
  wire n891_lo_buf_o2_n_spl_0;
  wire g722_n_spl_;
  wire g722_p_spl_;
  wire g726_p_spl_;
  wire n927_lo_buf_o2_p_spl_;
  wire n915_lo_buf_o2_p_spl_;
  wire n927_lo_buf_o2_n_spl_;
  wire n927_lo_buf_o2_n_spl_0;
  wire n915_lo_buf_o2_n_spl_;
  wire n915_lo_buf_o2_n_spl_0;
  wire g730_n_spl_;
  wire g730_p_spl_;
  wire n951_lo_buf_o2_p_spl_;
  wire n939_lo_buf_o2_p_spl_;
  wire n951_lo_buf_o2_n_spl_;
  wire n951_lo_buf_o2_n_spl_0;
  wire n939_lo_buf_o2_n_spl_;
  wire n939_lo_buf_o2_n_spl_0;
  wire g734_n_spl_;
  wire g734_p_spl_;
  wire g738_p_spl_;
  wire n975_lo_buf_o2_p_spl_;
  wire n963_lo_buf_o2_p_spl_;
  wire n975_lo_buf_o2_n_spl_;
  wire n975_lo_buf_o2_n_spl_0;
  wire n963_lo_buf_o2_n_spl_;
  wire n963_lo_buf_o2_n_spl_0;
  wire g742_n_spl_;
  wire g742_p_spl_;
  wire n999_lo_buf_o2_p_spl_;
  wire n987_lo_buf_o2_p_spl_;
  wire n999_lo_buf_o2_n_spl_;
  wire n999_lo_buf_o2_n_spl_0;
  wire n987_lo_buf_o2_n_spl_;
  wire n987_lo_buf_o2_n_spl_0;
  wire g746_n_spl_;
  wire g746_p_spl_;
  wire g750_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    n630_lo_p,
    n630_lo
  );


  not

  (
    n630_lo_n,
    n630_lo
  );


  buf

  (
    n642_lo_p,
    n642_lo
  );


  not

  (
    n642_lo_n,
    n642_lo
  );


  buf

  (
    n654_lo_p,
    n654_lo
  );


  not

  (
    n654_lo_n,
    n654_lo
  );


  buf

  (
    n666_lo_p,
    n666_lo
  );


  not

  (
    n666_lo_n,
    n666_lo
  );


  buf

  (
    n678_lo_p,
    n678_lo
  );


  not

  (
    n678_lo_n,
    n678_lo
  );


  buf

  (
    n690_lo_p,
    n690_lo
  );


  not

  (
    n690_lo_n,
    n690_lo
  );


  buf

  (
    n702_lo_p,
    n702_lo
  );


  not

  (
    n702_lo_n,
    n702_lo
  );


  buf

  (
    n714_lo_p,
    n714_lo
  );


  not

  (
    n714_lo_n,
    n714_lo
  );


  buf

  (
    n726_lo_p,
    n726_lo
  );


  not

  (
    n726_lo_n,
    n726_lo
  );


  buf

  (
    n738_lo_p,
    n738_lo
  );


  not

  (
    n738_lo_n,
    n738_lo
  );


  buf

  (
    n750_lo_p,
    n750_lo
  );


  not

  (
    n750_lo_n,
    n750_lo
  );


  buf

  (
    n762_lo_p,
    n762_lo
  );


  not

  (
    n762_lo_n,
    n762_lo
  );


  buf

  (
    n774_lo_p,
    n774_lo
  );


  not

  (
    n774_lo_n,
    n774_lo
  );


  buf

  (
    n786_lo_p,
    n786_lo
  );


  not

  (
    n786_lo_n,
    n786_lo
  );


  buf

  (
    n798_lo_p,
    n798_lo
  );


  not

  (
    n798_lo_n,
    n798_lo
  );


  buf

  (
    n810_lo_p,
    n810_lo
  );


  not

  (
    n810_lo_n,
    n810_lo
  );


  buf

  (
    n822_lo_p,
    n822_lo
  );


  not

  (
    n822_lo_n,
    n822_lo
  );


  buf

  (
    n834_lo_p,
    n834_lo
  );


  not

  (
    n834_lo_n,
    n834_lo
  );


  buf

  (
    n846_lo_p,
    n846_lo
  );


  not

  (
    n846_lo_n,
    n846_lo
  );


  buf

  (
    n858_lo_p,
    n858_lo
  );


  not

  (
    n858_lo_n,
    n858_lo
  );


  buf

  (
    n870_lo_p,
    n870_lo
  );


  not

  (
    n870_lo_n,
    n870_lo
  );


  buf

  (
    n882_lo_p,
    n882_lo
  );


  not

  (
    n882_lo_n,
    n882_lo
  );


  buf

  (
    n894_lo_p,
    n894_lo
  );


  not

  (
    n894_lo_n,
    n894_lo
  );


  buf

  (
    n906_lo_p,
    n906_lo
  );


  not

  (
    n906_lo_n,
    n906_lo
  );


  buf

  (
    n918_lo_p,
    n918_lo
  );


  not

  (
    n918_lo_n,
    n918_lo
  );


  buf

  (
    n930_lo_p,
    n930_lo
  );


  not

  (
    n930_lo_n,
    n930_lo
  );


  buf

  (
    n942_lo_p,
    n942_lo
  );


  not

  (
    n942_lo_n,
    n942_lo
  );


  buf

  (
    n954_lo_p,
    n954_lo
  );


  not

  (
    n954_lo_n,
    n954_lo
  );


  buf

  (
    n966_lo_p,
    n966_lo
  );


  not

  (
    n966_lo_n,
    n966_lo
  );


  buf

  (
    n978_lo_p,
    n978_lo
  );


  not

  (
    n978_lo_n,
    n978_lo
  );


  buf

  (
    n990_lo_p,
    n990_lo
  );


  not

  (
    n990_lo_n,
    n990_lo
  );


  buf

  (
    n1002_lo_p,
    n1002_lo
  );


  not

  (
    n1002_lo_n,
    n1002_lo
  );


  buf

  (
    n1005_lo_p,
    n1005_lo
  );


  not

  (
    n1005_lo_n,
    n1005_lo
  );


  buf

  (
    n1008_lo_p,
    n1008_lo
  );


  not

  (
    n1008_lo_n,
    n1008_lo
  );


  buf

  (
    n1017_lo_p,
    n1017_lo
  );


  not

  (
    n1017_lo_n,
    n1017_lo
  );


  buf

  (
    n1020_lo_p,
    n1020_lo
  );


  not

  (
    n1020_lo_n,
    n1020_lo
  );


  buf

  (
    n1029_lo_p,
    n1029_lo
  );


  not

  (
    n1029_lo_n,
    n1029_lo
  );


  buf

  (
    n1032_lo_p,
    n1032_lo
  );


  not

  (
    n1032_lo_n,
    n1032_lo
  );


  buf

  (
    n1041_lo_p,
    n1041_lo
  );


  not

  (
    n1041_lo_n,
    n1041_lo
  );


  buf

  (
    n1044_lo_p,
    n1044_lo
  );


  not

  (
    n1044_lo_n,
    n1044_lo
  );


  buf

  (
    n1053_lo_p,
    n1053_lo
  );


  not

  (
    n1053_lo_n,
    n1053_lo
  );


  buf

  (
    n1056_lo_p,
    n1056_lo
  );


  not

  (
    n1056_lo_n,
    n1056_lo
  );


  buf

  (
    n1065_lo_p,
    n1065_lo
  );


  not

  (
    n1065_lo_n,
    n1065_lo
  );


  buf

  (
    n1068_lo_p,
    n1068_lo
  );


  not

  (
    n1068_lo_n,
    n1068_lo
  );


  buf

  (
    n1077_lo_p,
    n1077_lo
  );


  not

  (
    n1077_lo_n,
    n1077_lo
  );


  buf

  (
    n1080_lo_p,
    n1080_lo
  );


  not

  (
    n1080_lo_n,
    n1080_lo
  );


  buf

  (
    n1089_lo_p,
    n1089_lo
  );


  not

  (
    n1089_lo_n,
    n1089_lo
  );


  buf

  (
    n1092_lo_p,
    n1092_lo
  );


  not

  (
    n1092_lo_n,
    n1092_lo
  );


  buf

  (
    n1101_lo_p,
    n1101_lo
  );


  not

  (
    n1101_lo_n,
    n1101_lo
  );


  buf

  (
    n1104_lo_p,
    n1104_lo
  );


  not

  (
    n1104_lo_n,
    n1104_lo
  );


  buf

  (
    n1837_o2_p,
    n1837_o2
  );


  not

  (
    n1837_o2_n,
    n1837_o2
  );


  buf

  (
    n1838_o2_p,
    n1838_o2
  );


  not

  (
    n1838_o2_n,
    n1838_o2
  );


  buf

  (
    n1839_o2_p,
    n1839_o2
  );


  not

  (
    n1839_o2_n,
    n1839_o2
  );


  buf

  (
    n1840_o2_p,
    n1840_o2
  );


  not

  (
    n1840_o2_n,
    n1840_o2
  );


  buf

  (
    n1841_o2_p,
    n1841_o2
  );


  not

  (
    n1841_o2_n,
    n1841_o2
  );


  buf

  (
    n1842_o2_p,
    n1842_o2
  );


  not

  (
    n1842_o2_n,
    n1842_o2
  );


  buf

  (
    n1843_o2_p,
    n1843_o2
  );


  not

  (
    n1843_o2_n,
    n1843_o2
  );


  buf

  (
    n1844_o2_p,
    n1844_o2
  );


  not

  (
    n1844_o2_n,
    n1844_o2
  );


  buf

  (
    n1845_o2_p,
    n1845_o2
  );


  not

  (
    n1845_o2_n,
    n1845_o2
  );


  buf

  (
    n1846_o2_p,
    n1846_o2
  );


  not

  (
    n1846_o2_n,
    n1846_o2
  );


  buf

  (
    n1847_o2_p,
    n1847_o2
  );


  not

  (
    n1847_o2_n,
    n1847_o2
  );


  buf

  (
    n1848_o2_p,
    n1848_o2
  );


  not

  (
    n1848_o2_n,
    n1848_o2
  );


  buf

  (
    n1849_o2_p,
    n1849_o2
  );


  not

  (
    n1849_o2_n,
    n1849_o2
  );


  buf

  (
    n1850_o2_p,
    n1850_o2
  );


  not

  (
    n1850_o2_n,
    n1850_o2
  );


  buf

  (
    n1851_o2_p,
    n1851_o2
  );


  not

  (
    n1851_o2_n,
    n1851_o2
  );


  buf

  (
    n1852_o2_p,
    n1852_o2
  );


  not

  (
    n1852_o2_n,
    n1852_o2
  );


  buf

  (
    n1853_o2_p,
    n1853_o2
  );


  not

  (
    n1853_o2_n,
    n1853_o2
  );


  buf

  (
    n1854_o2_p,
    n1854_o2
  );


  not

  (
    n1854_o2_n,
    n1854_o2
  );


  buf

  (
    n1855_o2_p,
    n1855_o2
  );


  not

  (
    n1855_o2_n,
    n1855_o2
  );


  buf

  (
    n1856_o2_p,
    n1856_o2
  );


  not

  (
    n1856_o2_n,
    n1856_o2
  );


  buf

  (
    n1857_o2_p,
    n1857_o2
  );


  not

  (
    n1857_o2_n,
    n1857_o2
  );


  buf

  (
    n1858_o2_p,
    n1858_o2
  );


  not

  (
    n1858_o2_n,
    n1858_o2
  );


  buf

  (
    n1859_o2_p,
    n1859_o2
  );


  not

  (
    n1859_o2_n,
    n1859_o2
  );


  buf

  (
    n1860_o2_p,
    n1860_o2
  );


  not

  (
    n1860_o2_n,
    n1860_o2
  );


  buf

  (
    n1861_o2_p,
    n1861_o2
  );


  not

  (
    n1861_o2_n,
    n1861_o2
  );


  buf

  (
    n1862_o2_p,
    n1862_o2
  );


  not

  (
    n1862_o2_n,
    n1862_o2
  );


  buf

  (
    n1863_o2_p,
    n1863_o2
  );


  not

  (
    n1863_o2_n,
    n1863_o2
  );


  buf

  (
    n1864_o2_p,
    n1864_o2
  );


  not

  (
    n1864_o2_n,
    n1864_o2
  );


  buf

  (
    n1865_o2_p,
    n1865_o2
  );


  not

  (
    n1865_o2_n,
    n1865_o2
  );


  buf

  (
    n1866_o2_p,
    n1866_o2
  );


  not

  (
    n1866_o2_n,
    n1866_o2
  );


  buf

  (
    n1867_o2_p,
    n1867_o2
  );


  not

  (
    n1867_o2_n,
    n1867_o2
  );


  buf

  (
    n1868_o2_p,
    n1868_o2
  );


  not

  (
    n1868_o2_n,
    n1868_o2
  );


  buf

  (
    G834_o2_p,
    G834_o2
  );


  not

  (
    G834_o2_n,
    G834_o2
  );


  buf

  (
    G847_o2_p,
    G847_o2
  );


  not

  (
    G847_o2_n,
    G847_o2
  );


  buf

  (
    G860_o2_p,
    G860_o2
  );


  not

  (
    G860_o2_n,
    G860_o2
  );


  buf

  (
    G873_o2_p,
    G873_o2
  );


  not

  (
    G873_o2_n,
    G873_o2
  );


  buf

  (
    G925_o2_p,
    G925_o2
  );


  not

  (
    G925_o2_n,
    G925_o2
  );


  buf

  (
    G886_o2_p,
    G886_o2
  );


  not

  (
    G886_o2_n,
    G886_o2
  );


  buf

  (
    G912_o2_p,
    G912_o2
  );


  not

  (
    G912_o2_n,
    G912_o2
  );


  buf

  (
    G899_o2_p,
    G899_o2
  );


  not

  (
    G899_o2_n,
    G899_o2
  );


  buf

  (
    n2151_o2_p,
    n2151_o2
  );


  not

  (
    n2151_o2_n,
    n2151_o2
  );


  buf

  (
    n2152_o2_p,
    n2152_o2
  );


  not

  (
    n2152_o2_n,
    n2152_o2
  );


  buf

  (
    n2153_o2_p,
    n2153_o2
  );


  not

  (
    n2153_o2_n,
    n2153_o2
  );


  buf

  (
    n2154_o2_p,
    n2154_o2
  );


  not

  (
    n2154_o2_n,
    n2154_o2
  );


  buf

  (
    n2155_o2_p,
    n2155_o2
  );


  not

  (
    n2155_o2_n,
    n2155_o2
  );


  buf

  (
    n2156_o2_p,
    n2156_o2
  );


  not

  (
    n2156_o2_n,
    n2156_o2
  );


  buf

  (
    n2157_o2_p,
    n2157_o2
  );


  not

  (
    n2157_o2_n,
    n2157_o2
  );


  buf

  (
    n2158_o2_p,
    n2158_o2
  );


  not

  (
    n2158_o2_n,
    n2158_o2
  );


  buf

  (
    n2159_o2_p,
    n2159_o2
  );


  not

  (
    n2159_o2_n,
    n2159_o2
  );


  buf

  (
    n2160_o2_p,
    n2160_o2
  );


  not

  (
    n2160_o2_n,
    n2160_o2
  );


  buf

  (
    n2161_o2_p,
    n2161_o2
  );


  not

  (
    n2161_o2_n,
    n2161_o2
  );


  buf

  (
    n2162_o2_p,
    n2162_o2
  );


  not

  (
    n2162_o2_n,
    n2162_o2
  );


  buf

  (
    n2163_o2_p,
    n2163_o2
  );


  not

  (
    n2163_o2_n,
    n2163_o2
  );


  buf

  (
    n2164_o2_p,
    n2164_o2
  );


  not

  (
    n2164_o2_n,
    n2164_o2
  );


  buf

  (
    n2165_o2_p,
    n2165_o2
  );


  not

  (
    n2165_o2_n,
    n2165_o2
  );


  buf

  (
    n2166_o2_p,
    n2166_o2
  );


  not

  (
    n2166_o2_n,
    n2166_o2
  );


  buf

  (
    n2167_o2_p,
    n2167_o2
  );


  not

  (
    n2167_o2_n,
    n2167_o2
  );


  buf

  (
    n2168_o2_p,
    n2168_o2
  );


  not

  (
    n2168_o2_n,
    n2168_o2
  );


  buf

  (
    n2169_o2_p,
    n2169_o2
  );


  not

  (
    n2169_o2_n,
    n2169_o2
  );


  buf

  (
    n2170_o2_p,
    n2170_o2
  );


  not

  (
    n2170_o2_n,
    n2170_o2
  );


  buf

  (
    n2171_o2_p,
    n2171_o2
  );


  not

  (
    n2171_o2_n,
    n2171_o2
  );


  buf

  (
    n2172_o2_p,
    n2172_o2
  );


  not

  (
    n2172_o2_n,
    n2172_o2
  );


  buf

  (
    n2173_o2_p,
    n2173_o2
  );


  not

  (
    n2173_o2_n,
    n2173_o2
  );


  buf

  (
    n2174_o2_p,
    n2174_o2
  );


  not

  (
    n2174_o2_n,
    n2174_o2
  );


  buf

  (
    n2175_o2_p,
    n2175_o2
  );


  not

  (
    n2175_o2_n,
    n2175_o2
  );


  buf

  (
    n2176_o2_p,
    n2176_o2
  );


  not

  (
    n2176_o2_n,
    n2176_o2
  );


  buf

  (
    n2177_o2_p,
    n2177_o2
  );


  not

  (
    n2177_o2_n,
    n2177_o2
  );


  buf

  (
    n2178_o2_p,
    n2178_o2
  );


  not

  (
    n2178_o2_n,
    n2178_o2
  );


  buf

  (
    n2179_o2_p,
    n2179_o2
  );


  not

  (
    n2179_o2_n,
    n2179_o2
  );


  buf

  (
    n2180_o2_p,
    n2180_o2
  );


  not

  (
    n2180_o2_n,
    n2180_o2
  );


  buf

  (
    n2181_o2_p,
    n2181_o2
  );


  not

  (
    n2181_o2_n,
    n2181_o2
  );


  buf

  (
    n2182_o2_p,
    n2182_o2
  );


  not

  (
    n2182_o2_n,
    n2182_o2
  );


  buf

  (
    G974_o2_p,
    G974_o2
  );


  not

  (
    G974_o2_n,
    G974_o2
  );


  buf

  (
    G976_o2_p,
    G976_o2
  );


  not

  (
    G976_o2_n,
    G976_o2
  );


  buf

  (
    G970_o2_p,
    G970_o2
  );


  not

  (
    G970_o2_n,
    G970_o2
  );


  buf

  (
    G972_o2_p,
    G972_o2
  );


  not

  (
    G972_o2_n,
    G972_o2
  );


  buf

  (
    G973_o2_p,
    G973_o2
  );


  not

  (
    G973_o2_n,
    G973_o2
  );


  buf

  (
    G977_o2_p,
    G977_o2
  );


  not

  (
    G977_o2_n,
    G977_o2
  );


  buf

  (
    G971_o2_p,
    G971_o2
  );


  not

  (
    G971_o2_n,
    G971_o2
  );


  buf

  (
    G975_o2_p,
    G975_o2
  );


  not

  (
    G975_o2_n,
    G975_o2
  );


  buf

  (
    G954_o2_p,
    G954_o2
  );


  not

  (
    G954_o2_n,
    G954_o2
  );


  buf

  (
    G956_o2_p,
    G956_o2
  );


  not

  (
    G956_o2_n,
    G956_o2
  );


  buf

  (
    G950_o2_p,
    G950_o2
  );


  not

  (
    G950_o2_n,
    G950_o2
  );


  buf

  (
    G952_o2_p,
    G952_o2
  );


  not

  (
    G952_o2_n,
    G952_o2
  );


  buf

  (
    G953_o2_p,
    G953_o2
  );


  not

  (
    G953_o2_n,
    G953_o2
  );


  buf

  (
    G957_o2_p,
    G957_o2
  );


  not

  (
    G957_o2_n,
    G957_o2
  );


  buf

  (
    G951_o2_p,
    G951_o2
  );


  not

  (
    G951_o2_n,
    G951_o2
  );


  buf

  (
    G955_o2_p,
    G955_o2
  );


  not

  (
    G955_o2_n,
    G955_o2
  );


  buf

  (
    G986_o2_p,
    G986_o2
  );


  not

  (
    G986_o2_n,
    G986_o2
  );


  buf

  (
    G991_o2_p,
    G991_o2
  );


  not

  (
    G991_o2_n,
    G991_o2
  );


  buf

  (
    G770_o2_p,
    G770_o2
  );


  not

  (
    G770_o2_n,
    G770_o2
  );


  buf

  (
    G773_o2_p,
    G773_o2
  );


  not

  (
    G773_o2_n,
    G773_o2
  );


  buf

  (
    G776_o2_p,
    G776_o2
  );


  not

  (
    G776_o2_n,
    G776_o2
  );


  buf

  (
    G779_o2_p,
    G779_o2
  );


  not

  (
    G779_o2_n,
    G779_o2
  );


  buf

  (
    G782_o2_p,
    G782_o2
  );


  not

  (
    G782_o2_n,
    G782_o2
  );


  buf

  (
    G785_o2_p,
    G785_o2
  );


  not

  (
    G785_o2_n,
    G785_o2
  );


  buf

  (
    G788_o2_p,
    G788_o2
  );


  not

  (
    G788_o2_n,
    G788_o2
  );


  buf

  (
    G791_o2_p,
    G791_o2
  );


  not

  (
    G791_o2_n,
    G791_o2
  );


  buf

  (
    G642_o2_p,
    G642_o2
  );


  not

  (
    G642_o2_n,
    G642_o2
  );


  buf

  (
    G645_o2_p,
    G645_o2
  );


  not

  (
    G645_o2_n,
    G645_o2
  );


  buf

  (
    G648_o2_p,
    G648_o2
  );


  not

  (
    G648_o2_n,
    G648_o2
  );


  buf

  (
    G651_o2_p,
    G651_o2
  );


  not

  (
    G651_o2_n,
    G651_o2
  );


  buf

  (
    G654_o2_p,
    G654_o2
  );


  not

  (
    G654_o2_n,
    G654_o2
  );


  buf

  (
    G657_o2_p,
    G657_o2
  );


  not

  (
    G657_o2_n,
    G657_o2
  );


  buf

  (
    G660_o2_p,
    G660_o2
  );


  not

  (
    G660_o2_n,
    G660_o2
  );


  buf

  (
    G663_o2_p,
    G663_o2
  );


  not

  (
    G663_o2_n,
    G663_o2
  );


  buf

  (
    G602_o2_p,
    G602_o2
  );


  not

  (
    G602_o2_n,
    G602_o2
  );


  buf

  (
    G607_o2_p,
    G607_o2
  );


  not

  (
    G607_o2_n,
    G607_o2
  );


  buf

  (
    G612_o2_p,
    G612_o2
  );


  not

  (
    G612_o2_n,
    G612_o2
  );


  buf

  (
    G617_o2_p,
    G617_o2
  );


  not

  (
    G617_o2_n,
    G617_o2
  );


  buf

  (
    G622_o2_p,
    G622_o2
  );


  not

  (
    G622_o2_n,
    G622_o2
  );


  buf

  (
    G627_o2_p,
    G627_o2
  );


  not

  (
    G627_o2_n,
    G627_o2
  );


  buf

  (
    G632_o2_p,
    G632_o2
  );


  not

  (
    G632_o2_n,
    G632_o2
  );


  buf

  (
    G637_o2_p,
    G637_o2
  );


  not

  (
    G637_o2_n,
    G637_o2
  );


  buf

  (
    n627_lo_buf_o2_p,
    n627_lo_buf_o2
  );


  not

  (
    n627_lo_buf_o2_n,
    n627_lo_buf_o2
  );


  buf

  (
    n639_lo_buf_o2_p,
    n639_lo_buf_o2
  );


  not

  (
    n639_lo_buf_o2_n,
    n639_lo_buf_o2
  );


  buf

  (
    n651_lo_buf_o2_p,
    n651_lo_buf_o2
  );


  not

  (
    n651_lo_buf_o2_n,
    n651_lo_buf_o2
  );


  buf

  (
    n663_lo_buf_o2_p,
    n663_lo_buf_o2
  );


  not

  (
    n663_lo_buf_o2_n,
    n663_lo_buf_o2
  );


  buf

  (
    n675_lo_buf_o2_p,
    n675_lo_buf_o2
  );


  not

  (
    n675_lo_buf_o2_n,
    n675_lo_buf_o2
  );


  buf

  (
    n687_lo_buf_o2_p,
    n687_lo_buf_o2
  );


  not

  (
    n687_lo_buf_o2_n,
    n687_lo_buf_o2
  );


  buf

  (
    n699_lo_buf_o2_p,
    n699_lo_buf_o2
  );


  not

  (
    n699_lo_buf_o2_n,
    n699_lo_buf_o2
  );


  buf

  (
    n711_lo_buf_o2_p,
    n711_lo_buf_o2
  );


  not

  (
    n711_lo_buf_o2_n,
    n711_lo_buf_o2
  );


  buf

  (
    n723_lo_buf_o2_p,
    n723_lo_buf_o2
  );


  not

  (
    n723_lo_buf_o2_n,
    n723_lo_buf_o2
  );


  buf

  (
    n735_lo_buf_o2_p,
    n735_lo_buf_o2
  );


  not

  (
    n735_lo_buf_o2_n,
    n735_lo_buf_o2
  );


  buf

  (
    n747_lo_buf_o2_p,
    n747_lo_buf_o2
  );


  not

  (
    n747_lo_buf_o2_n,
    n747_lo_buf_o2
  );


  buf

  (
    n759_lo_buf_o2_p,
    n759_lo_buf_o2
  );


  not

  (
    n759_lo_buf_o2_n,
    n759_lo_buf_o2
  );


  buf

  (
    n771_lo_buf_o2_p,
    n771_lo_buf_o2
  );


  not

  (
    n771_lo_buf_o2_n,
    n771_lo_buf_o2
  );


  buf

  (
    n783_lo_buf_o2_p,
    n783_lo_buf_o2
  );


  not

  (
    n783_lo_buf_o2_n,
    n783_lo_buf_o2
  );


  buf

  (
    n795_lo_buf_o2_p,
    n795_lo_buf_o2
  );


  not

  (
    n795_lo_buf_o2_n,
    n795_lo_buf_o2
  );


  buf

  (
    n807_lo_buf_o2_p,
    n807_lo_buf_o2
  );


  not

  (
    n807_lo_buf_o2_n,
    n807_lo_buf_o2
  );


  buf

  (
    n819_lo_buf_o2_p,
    n819_lo_buf_o2
  );


  not

  (
    n819_lo_buf_o2_n,
    n819_lo_buf_o2
  );


  buf

  (
    n831_lo_buf_o2_p,
    n831_lo_buf_o2
  );


  not

  (
    n831_lo_buf_o2_n,
    n831_lo_buf_o2
  );


  buf

  (
    n843_lo_buf_o2_p,
    n843_lo_buf_o2
  );


  not

  (
    n843_lo_buf_o2_n,
    n843_lo_buf_o2
  );


  buf

  (
    n855_lo_buf_o2_p,
    n855_lo_buf_o2
  );


  not

  (
    n855_lo_buf_o2_n,
    n855_lo_buf_o2
  );


  buf

  (
    n867_lo_buf_o2_p,
    n867_lo_buf_o2
  );


  not

  (
    n867_lo_buf_o2_n,
    n867_lo_buf_o2
  );


  buf

  (
    n879_lo_buf_o2_p,
    n879_lo_buf_o2
  );


  not

  (
    n879_lo_buf_o2_n,
    n879_lo_buf_o2
  );


  buf

  (
    n891_lo_buf_o2_p,
    n891_lo_buf_o2
  );


  not

  (
    n891_lo_buf_o2_n,
    n891_lo_buf_o2
  );


  buf

  (
    n903_lo_buf_o2_p,
    n903_lo_buf_o2
  );


  not

  (
    n903_lo_buf_o2_n,
    n903_lo_buf_o2
  );


  buf

  (
    n915_lo_buf_o2_p,
    n915_lo_buf_o2
  );


  not

  (
    n915_lo_buf_o2_n,
    n915_lo_buf_o2
  );


  buf

  (
    n927_lo_buf_o2_p,
    n927_lo_buf_o2
  );


  not

  (
    n927_lo_buf_o2_n,
    n927_lo_buf_o2
  );


  buf

  (
    n939_lo_buf_o2_p,
    n939_lo_buf_o2
  );


  not

  (
    n939_lo_buf_o2_n,
    n939_lo_buf_o2
  );


  buf

  (
    n951_lo_buf_o2_p,
    n951_lo_buf_o2
  );


  not

  (
    n951_lo_buf_o2_n,
    n951_lo_buf_o2
  );


  buf

  (
    n963_lo_buf_o2_p,
    n963_lo_buf_o2
  );


  not

  (
    n963_lo_buf_o2_n,
    n963_lo_buf_o2
  );


  buf

  (
    n975_lo_buf_o2_p,
    n975_lo_buf_o2
  );


  not

  (
    n975_lo_buf_o2_n,
    n975_lo_buf_o2
  );


  buf

  (
    n987_lo_buf_o2_p,
    n987_lo_buf_o2
  );


  not

  (
    n987_lo_buf_o2_n,
    n987_lo_buf_o2
  );


  buf

  (
    n999_lo_buf_o2_p,
    n999_lo_buf_o2
  );


  not

  (
    n999_lo_buf_o2_n,
    n999_lo_buf_o2
  );


  and

  (
    g238_p,
    G950_o2_n,
    G925_o2_p_spl_00
  );


  or

  (
    g238_n,
    G950_o2_p,
    G925_o2_n_spl_00
  );


  and

  (
    g239_p,
    g238_p,
    G912_o2_p_spl_00
  );


  or

  (
    g239_n,
    g238_n,
    G912_o2_n_spl_00
  );


  and

  (
    g240_p,
    g239_p,
    G951_o2_n
  );


  or

  (
    g240_n,
    g239_n,
    G951_o2_p
  );


  and

  (
    g241_p,
    g240_p,
    G986_o2_p_spl_0
  );


  or

  (
    g241_n,
    g240_n,
    G986_o2_n_spl_0
  );


  and

  (
    g242_p,
    g241_p_spl_0,
    G834_o2_p_spl_00
  );


  or

  (
    g242_n,
    g241_n_spl_0,
    G834_o2_n_spl_00
  );


  or

  (
    g243_n,
    g242_n,
    n630_lo_n
  );


  and

  (
    g244_p,
    g243_n_spl_,
    n630_lo_p
  );


  and

  (
    g245_p,
    g243_n_spl_,
    g242_p
  );


  or

  (
    g246_n,
    g245_p,
    g244_p
  );


  and

  (
    g247_p,
    g241_p_spl_0,
    G847_o2_p_spl_00
  );


  or

  (
    g247_n,
    g241_n_spl_0,
    G847_o2_n_spl_00
  );


  or

  (
    g248_n,
    g247_n,
    n642_lo_n
  );


  and

  (
    g249_p,
    g248_n_spl_,
    n642_lo_p
  );


  and

  (
    g250_p,
    g248_n_spl_,
    g247_p
  );


  or

  (
    g251_n,
    g250_p,
    g249_p
  );


  and

  (
    g252_p,
    g241_p_spl_1,
    G860_o2_p_spl_00
  );


  or

  (
    g252_n,
    g241_n_spl_1,
    G860_o2_n_spl_00
  );


  or

  (
    g253_n,
    g252_n,
    n654_lo_n
  );


  and

  (
    g254_p,
    g253_n_spl_,
    n654_lo_p
  );


  and

  (
    g255_p,
    g253_n_spl_,
    g252_p
  );


  or

  (
    g256_n,
    g255_p,
    g254_p
  );


  and

  (
    g257_p,
    g241_p_spl_1,
    G873_o2_p_spl_00
  );


  or

  (
    g257_n,
    g241_n_spl_1,
    G873_o2_n_spl_00
  );


  or

  (
    g258_n,
    g257_n,
    n666_lo_n
  );


  and

  (
    g259_p,
    g258_n_spl_,
    n666_lo_p
  );


  and

  (
    g260_p,
    g258_n_spl_,
    g257_p
  );


  or

  (
    g261_n,
    g260_p,
    g259_p
  );


  and

  (
    g262_p,
    G952_o2_n,
    G925_o2_p_spl_00
  );


  or

  (
    g262_n,
    G952_o2_p,
    G925_o2_n_spl_00
  );


  and

  (
    g263_p,
    g262_p,
    G953_o2_n
  );


  or

  (
    g263_n,
    g262_n,
    G953_o2_p
  );


  and

  (
    g264_p,
    g263_p,
    G899_o2_p_spl_00
  );


  or

  (
    g264_n,
    g263_n,
    G899_o2_n_spl_00
  );


  and

  (
    g265_p,
    g264_p,
    G986_o2_p_spl_0
  );


  or

  (
    g265_n,
    g264_n,
    G986_o2_n_spl_0
  );


  and

  (
    g266_p,
    g265_p_spl_0,
    G834_o2_p_spl_00
  );


  or

  (
    g266_n,
    g265_n_spl_0,
    G834_o2_n_spl_00
  );


  or

  (
    g267_n,
    g266_n,
    n678_lo_n
  );


  and

  (
    g268_p,
    g267_n_spl_,
    n678_lo_p
  );


  and

  (
    g269_p,
    g267_n_spl_,
    g266_p
  );


  or

  (
    g270_n,
    g269_p,
    g268_p
  );


  and

  (
    g271_p,
    g265_p_spl_0,
    G847_o2_p_spl_00
  );


  or

  (
    g271_n,
    g265_n_spl_0,
    G847_o2_n_spl_00
  );


  or

  (
    g272_n,
    g271_n,
    n690_lo_n
  );


  and

  (
    g273_p,
    g272_n_spl_,
    n690_lo_p
  );


  and

  (
    g274_p,
    g272_n_spl_,
    g271_p
  );


  or

  (
    g275_n,
    g274_p,
    g273_p
  );


  and

  (
    g276_p,
    g265_p_spl_1,
    G860_o2_p_spl_00
  );


  or

  (
    g276_n,
    g265_n_spl_1,
    G860_o2_n_spl_00
  );


  or

  (
    g277_n,
    g276_n,
    n702_lo_n
  );


  and

  (
    g278_p,
    g277_n_spl_,
    n702_lo_p
  );


  and

  (
    g279_p,
    g277_n_spl_,
    g276_p
  );


  or

  (
    g280_n,
    g279_p,
    g278_p
  );


  and

  (
    g281_p,
    g265_p_spl_1,
    G873_o2_p_spl_00
  );


  or

  (
    g281_n,
    g265_n_spl_1,
    G873_o2_n_spl_00
  );


  or

  (
    g282_n,
    g281_n,
    n714_lo_n
  );


  and

  (
    g283_p,
    g282_n_spl_,
    n714_lo_p
  );


  and

  (
    g284_p,
    g282_n_spl_,
    g281_p
  );


  or

  (
    g285_n,
    g284_p,
    g283_p
  );


  and

  (
    g286_p,
    G954_o2_n,
    G886_o2_p_spl_00
  );


  or

  (
    g286_n,
    G954_o2_p,
    G886_o2_n_spl_00
  );


  and

  (
    g287_p,
    g286_p,
    G912_o2_p_spl_00
  );


  or

  (
    g287_n,
    g286_n,
    G912_o2_n_spl_00
  );


  and

  (
    g288_p,
    g287_p,
    G955_o2_n
  );


  or

  (
    g288_n,
    g287_n,
    G955_o2_p
  );


  and

  (
    g289_p,
    g288_p,
    G986_o2_p_spl_1
  );


  or

  (
    g289_n,
    g288_n,
    G986_o2_n_spl_1
  );


  and

  (
    g290_p,
    g289_p_spl_0,
    G834_o2_p_spl_01
  );


  or

  (
    g290_n,
    g289_n_spl_0,
    G834_o2_n_spl_01
  );


  or

  (
    g291_n,
    g290_n,
    n726_lo_n
  );


  and

  (
    g292_p,
    g291_n_spl_,
    n726_lo_p
  );


  and

  (
    g293_p,
    g291_n_spl_,
    g290_p
  );


  or

  (
    g294_n,
    g293_p,
    g292_p
  );


  and

  (
    g295_p,
    g289_p_spl_0,
    G847_o2_p_spl_01
  );


  or

  (
    g295_n,
    g289_n_spl_0,
    G847_o2_n_spl_01
  );


  or

  (
    g296_n,
    g295_n,
    n738_lo_n
  );


  and

  (
    g297_p,
    g296_n_spl_,
    n738_lo_p
  );


  and

  (
    g298_p,
    g296_n_spl_,
    g295_p
  );


  or

  (
    g299_n,
    g298_p,
    g297_p
  );


  and

  (
    g300_p,
    g289_p_spl_1,
    G860_o2_p_spl_01
  );


  or

  (
    g300_n,
    g289_n_spl_1,
    G860_o2_n_spl_01
  );


  or

  (
    g301_n,
    g300_n,
    n750_lo_n
  );


  and

  (
    g302_p,
    g301_n_spl_,
    n750_lo_p
  );


  and

  (
    g303_p,
    g301_n_spl_,
    g300_p
  );


  or

  (
    g304_n,
    g303_p,
    g302_p
  );


  and

  (
    g305_p,
    g289_p_spl_1,
    G873_o2_p_spl_01
  );


  or

  (
    g305_n,
    g289_n_spl_1,
    G873_o2_n_spl_01
  );


  or

  (
    g306_n,
    g305_n,
    n762_lo_n
  );


  and

  (
    g307_p,
    g306_n_spl_,
    n762_lo_p
  );


  and

  (
    g308_p,
    g306_n_spl_,
    g305_p
  );


  or

  (
    g309_n,
    g308_p,
    g307_p
  );


  and

  (
    g310_p,
    G956_o2_n,
    G886_o2_p_spl_00
  );


  or

  (
    g310_n,
    G956_o2_p,
    G886_o2_n_spl_00
  );


  and

  (
    g311_p,
    g310_p,
    G957_o2_n
  );


  or

  (
    g311_n,
    g310_n,
    G957_o2_p
  );


  and

  (
    g312_p,
    g311_p,
    G899_o2_p_spl_00
  );


  or

  (
    g312_n,
    g311_n,
    G899_o2_n_spl_00
  );


  and

  (
    g313_p,
    g312_p,
    G986_o2_p_spl_1
  );


  or

  (
    g313_n,
    g312_n,
    G986_o2_n_spl_1
  );


  and

  (
    g314_p,
    g313_p_spl_0,
    G834_o2_p_spl_01
  );


  or

  (
    g314_n,
    g313_n_spl_0,
    G834_o2_n_spl_01
  );


  or

  (
    g315_n,
    g314_n,
    n774_lo_n
  );


  and

  (
    g316_p,
    g315_n_spl_,
    n774_lo_p
  );


  and

  (
    g317_p,
    g315_n_spl_,
    g314_p
  );


  or

  (
    g318_n,
    g317_p,
    g316_p
  );


  and

  (
    g319_p,
    g313_p_spl_0,
    G847_o2_p_spl_01
  );


  or

  (
    g319_n,
    g313_n_spl_0,
    G847_o2_n_spl_01
  );


  or

  (
    g320_n,
    g319_n,
    n786_lo_n
  );


  and

  (
    g321_p,
    g320_n_spl_,
    n786_lo_p
  );


  and

  (
    g322_p,
    g320_n_spl_,
    g319_p
  );


  or

  (
    g323_n,
    g322_p,
    g321_p
  );


  and

  (
    g324_p,
    g313_p_spl_1,
    G860_o2_p_spl_01
  );


  or

  (
    g324_n,
    g313_n_spl_1,
    G860_o2_n_spl_01
  );


  or

  (
    g325_n,
    g324_n,
    n798_lo_n
  );


  and

  (
    g326_p,
    g325_n_spl_,
    n798_lo_p
  );


  and

  (
    g327_p,
    g325_n_spl_,
    g324_p
  );


  or

  (
    g328_n,
    g327_p,
    g326_p
  );


  and

  (
    g329_p,
    g313_p_spl_1,
    G873_o2_p_spl_01
  );


  or

  (
    g329_n,
    g313_n_spl_1,
    G873_o2_n_spl_01
  );


  or

  (
    g330_n,
    g329_n,
    n810_lo_n
  );


  and

  (
    g331_p,
    g330_n_spl_,
    n810_lo_p
  );


  and

  (
    g332_p,
    g330_n_spl_,
    g329_p
  );


  or

  (
    g333_n,
    g332_p,
    g331_p
  );


  and

  (
    g334_p,
    G970_o2_n,
    G834_o2_p_spl_1
  );


  or

  (
    g334_n,
    G970_o2_p,
    G834_o2_n_spl_1
  );


  and

  (
    g335_p,
    g334_p,
    G860_o2_p_spl_1
  );


  or

  (
    g335_n,
    g334_n,
    G860_o2_n_spl_1
  );


  and

  (
    g336_p,
    g335_p,
    G971_o2_n
  );


  or

  (
    g336_n,
    g335_n,
    G971_o2_p
  );


  and

  (
    g337_p,
    g336_p,
    G991_o2_p_spl_0
  );


  or

  (
    g337_n,
    g336_n,
    G991_o2_n_spl_0
  );


  and

  (
    g338_p,
    g337_p_spl_0,
    G925_o2_p_spl_01
  );


  or

  (
    g338_n,
    g337_n_spl_0,
    G925_o2_n_spl_01
  );


  or

  (
    g339_n,
    g338_n,
    n822_lo_n
  );


  and

  (
    g340_p,
    g339_n_spl_,
    n822_lo_p
  );


  and

  (
    g341_p,
    g339_n_spl_,
    g338_p
  );


  or

  (
    g342_n,
    g341_p,
    g340_p
  );


  and

  (
    g343_p,
    g337_p_spl_0,
    G886_o2_p_spl_01
  );


  or

  (
    g343_n,
    g337_n_spl_0,
    G886_o2_n_spl_01
  );


  or

  (
    g344_n,
    g343_n,
    n834_lo_n
  );


  and

  (
    g345_p,
    g344_n_spl_,
    n834_lo_p
  );


  and

  (
    g346_p,
    g344_n_spl_,
    g343_p
  );


  or

  (
    g347_n,
    g346_p,
    g345_p
  );


  and

  (
    g348_p,
    g337_p_spl_1,
    G912_o2_p_spl_01
  );


  or

  (
    g348_n,
    g337_n_spl_1,
    G912_o2_n_spl_01
  );


  or

  (
    g349_n,
    g348_n,
    n846_lo_n
  );


  and

  (
    g350_p,
    g349_n_spl_,
    n846_lo_p
  );


  and

  (
    g351_p,
    g349_n_spl_,
    g348_p
  );


  or

  (
    g352_n,
    g351_p,
    g350_p
  );


  and

  (
    g353_p,
    g337_p_spl_1,
    G899_o2_p_spl_01
  );


  or

  (
    g353_n,
    g337_n_spl_1,
    G899_o2_n_spl_01
  );


  or

  (
    g354_n,
    g353_n,
    n858_lo_n
  );


  and

  (
    g355_p,
    g354_n_spl_,
    n858_lo_p
  );


  and

  (
    g356_p,
    g354_n_spl_,
    g353_p
  );


  or

  (
    g357_n,
    g356_p,
    g355_p
  );


  and

  (
    g358_p,
    G972_o2_n,
    G834_o2_p_spl_1
  );


  or

  (
    g358_n,
    G972_o2_p,
    G834_o2_n_spl_1
  );


  and

  (
    g359_p,
    g358_p,
    G973_o2_n
  );


  or

  (
    g359_n,
    g358_n,
    G973_o2_p
  );


  and

  (
    g360_p,
    g359_p,
    G873_o2_p_spl_1
  );


  or

  (
    g360_n,
    g359_n,
    G873_o2_n_spl_1
  );


  and

  (
    g361_p,
    g360_p,
    G991_o2_p_spl_0
  );


  or

  (
    g361_n,
    g360_n,
    G991_o2_n_spl_0
  );


  and

  (
    g362_p,
    g361_p_spl_0,
    G925_o2_p_spl_01
  );


  or

  (
    g362_n,
    g361_n_spl_0,
    G925_o2_n_spl_01
  );


  or

  (
    g363_n,
    g362_n,
    n870_lo_n
  );


  and

  (
    g364_p,
    g363_n_spl_,
    n870_lo_p
  );


  and

  (
    g365_p,
    g363_n_spl_,
    g362_p
  );


  or

  (
    g366_n,
    g365_p,
    g364_p
  );


  and

  (
    g367_p,
    g361_p_spl_0,
    G886_o2_p_spl_01
  );


  or

  (
    g367_n,
    g361_n_spl_0,
    G886_o2_n_spl_01
  );


  or

  (
    g368_n,
    g367_n,
    n882_lo_n
  );


  and

  (
    g369_p,
    g368_n_spl_,
    n882_lo_p
  );


  and

  (
    g370_p,
    g368_n_spl_,
    g367_p
  );


  or

  (
    g371_n,
    g370_p,
    g369_p
  );


  and

  (
    g372_p,
    g361_p_spl_1,
    G912_o2_p_spl_01
  );


  or

  (
    g372_n,
    g361_n_spl_1,
    G912_o2_n_spl_01
  );


  or

  (
    g373_n,
    g372_n,
    n894_lo_n
  );


  and

  (
    g374_p,
    g373_n_spl_,
    n894_lo_p
  );


  and

  (
    g375_p,
    g373_n_spl_,
    g372_p
  );


  or

  (
    g376_n,
    g375_p,
    g374_p
  );


  and

  (
    g377_p,
    g361_p_spl_1,
    G899_o2_p_spl_01
  );


  or

  (
    g377_n,
    g361_n_spl_1,
    G899_o2_n_spl_01
  );


  or

  (
    g378_n,
    g377_n,
    n906_lo_n
  );


  and

  (
    g379_p,
    g378_n_spl_,
    n906_lo_p
  );


  and

  (
    g380_p,
    g378_n_spl_,
    g377_p
  );


  or

  (
    g381_n,
    g380_p,
    g379_p
  );


  and

  (
    g382_p,
    G974_o2_n,
    G847_o2_p_spl_1
  );


  or

  (
    g382_n,
    G974_o2_p,
    G847_o2_n_spl_1
  );


  and

  (
    g383_p,
    g382_p,
    G860_o2_p_spl_1
  );


  or

  (
    g383_n,
    g382_n,
    G860_o2_n_spl_1
  );


  and

  (
    g384_p,
    g383_p,
    G975_o2_n
  );


  or

  (
    g384_n,
    g383_n,
    G975_o2_p
  );


  and

  (
    g385_p,
    g384_p,
    G991_o2_p_spl_1
  );


  or

  (
    g385_n,
    g384_n,
    G991_o2_n_spl_1
  );


  and

  (
    g386_p,
    g385_p_spl_0,
    G925_o2_p_spl_1
  );


  or

  (
    g386_n,
    g385_n_spl_0,
    G925_o2_n_spl_1
  );


  or

  (
    g387_n,
    g386_n,
    n918_lo_n
  );


  and

  (
    g388_p,
    g387_n_spl_,
    n918_lo_p
  );


  and

  (
    g389_p,
    g387_n_spl_,
    g386_p
  );


  or

  (
    g390_n,
    g389_p,
    g388_p
  );


  and

  (
    g391_p,
    g385_p_spl_0,
    G886_o2_p_spl_1
  );


  or

  (
    g391_n,
    g385_n_spl_0,
    G886_o2_n_spl_1
  );


  or

  (
    g392_n,
    g391_n,
    n930_lo_n
  );


  and

  (
    g393_p,
    g392_n_spl_,
    n930_lo_p
  );


  and

  (
    g394_p,
    g392_n_spl_,
    g391_p
  );


  or

  (
    g395_n,
    g394_p,
    g393_p
  );


  and

  (
    g396_p,
    g385_p_spl_1,
    G912_o2_p_spl_1
  );


  or

  (
    g396_n,
    g385_n_spl_1,
    G912_o2_n_spl_1
  );


  or

  (
    g397_n,
    g396_n,
    n942_lo_n
  );


  and

  (
    g398_p,
    g397_n_spl_,
    n942_lo_p
  );


  and

  (
    g399_p,
    g397_n_spl_,
    g396_p
  );


  or

  (
    g400_n,
    g399_p,
    g398_p
  );


  and

  (
    g401_p,
    g385_p_spl_1,
    G899_o2_p_spl_1
  );


  or

  (
    g401_n,
    g385_n_spl_1,
    G899_o2_n_spl_1
  );


  or

  (
    g402_n,
    g401_n,
    n954_lo_n
  );


  and

  (
    g403_p,
    g402_n_spl_,
    n954_lo_p
  );


  and

  (
    g404_p,
    g402_n_spl_,
    g401_p
  );


  or

  (
    g405_n,
    g404_p,
    g403_p
  );


  and

  (
    g406_p,
    G976_o2_n,
    G847_o2_p_spl_1
  );


  or

  (
    g406_n,
    G976_o2_p,
    G847_o2_n_spl_1
  );


  and

  (
    g407_p,
    g406_p,
    G977_o2_n
  );


  or

  (
    g407_n,
    g406_n,
    G977_o2_p
  );


  and

  (
    g408_p,
    g407_p,
    G873_o2_p_spl_1
  );


  or

  (
    g408_n,
    g407_n,
    G873_o2_n_spl_1
  );


  and

  (
    g409_p,
    g408_p,
    G991_o2_p_spl_1
  );


  or

  (
    g409_n,
    g408_n,
    G991_o2_n_spl_1
  );


  and

  (
    g410_p,
    g409_p_spl_0,
    G925_o2_p_spl_1
  );


  or

  (
    g410_n,
    g409_n_spl_0,
    G925_o2_n_spl_1
  );


  or

  (
    g411_n,
    g410_n,
    n966_lo_n
  );


  and

  (
    g412_p,
    g411_n_spl_,
    n966_lo_p
  );


  and

  (
    g413_p,
    g411_n_spl_,
    g410_p
  );


  or

  (
    g414_n,
    g413_p,
    g412_p
  );


  and

  (
    g415_p,
    g409_p_spl_0,
    G886_o2_p_spl_1
  );


  or

  (
    g415_n,
    g409_n_spl_0,
    G886_o2_n_spl_1
  );


  or

  (
    g416_n,
    g415_n,
    n978_lo_n
  );


  and

  (
    g417_p,
    g416_n_spl_,
    n978_lo_p
  );


  and

  (
    g418_p,
    g416_n_spl_,
    g415_p
  );


  or

  (
    g419_n,
    g418_p,
    g417_p
  );


  and

  (
    g420_p,
    g409_p_spl_1,
    G912_o2_p_spl_1
  );


  or

  (
    g420_n,
    g409_n_spl_1,
    G912_o2_n_spl_1
  );


  or

  (
    g421_n,
    g420_n,
    n990_lo_n
  );


  and

  (
    g422_p,
    g421_n_spl_,
    n990_lo_p
  );


  and

  (
    g423_p,
    g421_n_spl_,
    g420_p
  );


  or

  (
    g424_n,
    g423_p,
    g422_p
  );


  and

  (
    g425_p,
    g409_p_spl_1,
    G899_o2_p_spl_1
  );


  or

  (
    g425_n,
    g409_n_spl_1,
    G899_o2_n_spl_1
  );


  or

  (
    g426_n,
    g425_n,
    n1002_lo_n
  );


  and

  (
    g427_p,
    g426_n_spl_,
    n1002_lo_p
  );


  and

  (
    g428_p,
    g426_n_spl_,
    g425_p
  );


  or

  (
    g429_n,
    g428_p,
    g427_p
  );


  and

  (
    g430_p,
    G642_o2_p_spl_,
    G770_o2_p_spl_
  );


  or

  (
    g430_n,
    G642_o2_n_spl_,
    G770_o2_n_spl_
  );


  and

  (
    g431_p,
    g430_n_spl_,
    G642_o2_p_spl_
  );


  or

  (
    g431_n,
    g430_p_spl_,
    G642_o2_n_spl_
  );


  and

  (
    g432_p,
    g430_n_spl_,
    G770_o2_p_spl_
  );


  or

  (
    g432_n,
    g430_p_spl_,
    G770_o2_n_spl_
  );


  and

  (
    g433_p,
    g432_n,
    g431_n
  );


  or

  (
    g433_n,
    g432_p,
    g431_p
  );


  and

  (
    g434_p,
    G645_o2_p_spl_,
    G773_o2_p_spl_
  );


  or

  (
    g434_n,
    G645_o2_n_spl_,
    G773_o2_n_spl_
  );


  and

  (
    g435_p,
    g434_n_spl_,
    G645_o2_p_spl_
  );


  or

  (
    g435_n,
    g434_p_spl_,
    G645_o2_n_spl_
  );


  and

  (
    g436_p,
    g434_n_spl_,
    G773_o2_p_spl_
  );


  or

  (
    g436_n,
    g434_p_spl_,
    G773_o2_n_spl_
  );


  and

  (
    g437_p,
    g436_n,
    g435_n
  );


  or

  (
    g437_n,
    g436_p,
    g435_p
  );


  and

  (
    g438_p,
    G648_o2_p_spl_,
    G776_o2_p_spl_
  );


  or

  (
    g438_n,
    G648_o2_n_spl_,
    G776_o2_n_spl_
  );


  and

  (
    g439_p,
    g438_n_spl_,
    G648_o2_p_spl_
  );


  or

  (
    g439_n,
    g438_p_spl_,
    G648_o2_n_spl_
  );


  and

  (
    g440_p,
    g438_n_spl_,
    G776_o2_p_spl_
  );


  or

  (
    g440_n,
    g438_p_spl_,
    G776_o2_n_spl_
  );


  and

  (
    g441_p,
    g440_n,
    g439_n
  );


  or

  (
    g441_n,
    g440_p,
    g439_p
  );


  and

  (
    g442_p,
    G651_o2_p_spl_,
    G779_o2_p_spl_
  );


  or

  (
    g442_n,
    G651_o2_n_spl_,
    G779_o2_n_spl_
  );


  and

  (
    g443_p,
    g442_n_spl_,
    G651_o2_p_spl_
  );


  or

  (
    g443_n,
    g442_p_spl_,
    G651_o2_n_spl_
  );


  and

  (
    g444_p,
    g442_n_spl_,
    G779_o2_p_spl_
  );


  or

  (
    g444_n,
    g442_p_spl_,
    G779_o2_n_spl_
  );


  and

  (
    g445_p,
    g444_n,
    g443_n
  );


  or

  (
    g445_n,
    g444_p,
    g443_p
  );


  and

  (
    g446_p,
    G654_o2_p_spl_,
    G782_o2_p_spl_
  );


  or

  (
    g446_n,
    G654_o2_n_spl_,
    G782_o2_n_spl_
  );


  and

  (
    g447_p,
    g446_n_spl_,
    G654_o2_p_spl_
  );


  or

  (
    g447_n,
    g446_p_spl_,
    G654_o2_n_spl_
  );


  and

  (
    g448_p,
    g446_n_spl_,
    G782_o2_p_spl_
  );


  or

  (
    g448_n,
    g446_p_spl_,
    G782_o2_n_spl_
  );


  and

  (
    g449_p,
    g448_n,
    g447_n
  );


  or

  (
    g449_n,
    g448_p,
    g447_p
  );


  and

  (
    g450_p,
    G657_o2_p_spl_,
    G785_o2_p_spl_
  );


  or

  (
    g450_n,
    G657_o2_n_spl_,
    G785_o2_n_spl_
  );


  and

  (
    g451_p,
    g450_n_spl_,
    G657_o2_p_spl_
  );


  or

  (
    g451_n,
    g450_p_spl_,
    G657_o2_n_spl_
  );


  and

  (
    g452_p,
    g450_n_spl_,
    G785_o2_p_spl_
  );


  or

  (
    g452_n,
    g450_p_spl_,
    G785_o2_n_spl_
  );


  and

  (
    g453_p,
    g452_n,
    g451_n
  );


  or

  (
    g453_n,
    g452_p,
    g451_p
  );


  and

  (
    g454_p,
    G660_o2_p_spl_,
    G788_o2_p_spl_
  );


  or

  (
    g454_n,
    G660_o2_n_spl_,
    G788_o2_n_spl_
  );


  and

  (
    g455_p,
    g454_n_spl_,
    G660_o2_p_spl_
  );


  or

  (
    g455_n,
    g454_p_spl_,
    G660_o2_n_spl_
  );


  and

  (
    g456_p,
    g454_n_spl_,
    G788_o2_p_spl_
  );


  or

  (
    g456_n,
    g454_p_spl_,
    G788_o2_n_spl_
  );


  and

  (
    g457_p,
    g456_n,
    g455_n
  );


  or

  (
    g457_n,
    g456_p,
    g455_p
  );


  and

  (
    g458_p,
    G663_o2_p_spl_,
    G791_o2_p_spl_
  );


  or

  (
    g458_n,
    G663_o2_n_spl_,
    G791_o2_n_spl_
  );


  and

  (
    g459_p,
    g458_n_spl_,
    G663_o2_p_spl_
  );


  or

  (
    g459_n,
    g458_p_spl_,
    G663_o2_n_spl_
  );


  and

  (
    g460_p,
    g458_n_spl_,
    G791_o2_p_spl_
  );


  or

  (
    g460_n,
    g458_p_spl_,
    G791_o2_n_spl_
  );


  and

  (
    g461_p,
    g460_n,
    g459_n
  );


  or

  (
    g461_n,
    g460_p,
    g459_p
  );


  or

  (
    g462_n,
    g437_n_spl_,
    g433_n_spl_
  );


  or

  (
    g463_n,
    g462_n_spl_,
    g441_n_spl_0
  );


  or

  (
    g464_n,
    g463_n,
    g445_p_spl_0
  );


  or

  (
    g465_n,
    g462_n_spl_,
    g441_p_spl_0
  );


  or

  (
    g466_n,
    g465_n,
    g445_n_spl_0
  );


  or

  (
    g467_n,
    g437_p_spl_0,
    g433_n_spl_
  );


  or

  (
    g468_n,
    g467_n,
    g441_n_spl_0
  );


  or

  (
    g469_n,
    g468_n,
    g445_n_spl_0
  );


  or

  (
    g470_n,
    g437_n_spl_,
    g433_p_spl_0
  );


  or

  (
    g471_n,
    g470_n,
    g441_n_spl_
  );


  or

  (
    g472_n,
    g471_n,
    g445_n_spl_
  );


  and

  (
    g473_p,
    g466_n,
    g464_n
  );


  and

  (
    g474_p,
    g473_p,
    g469_n
  );


  and

  (
    g475_p,
    g474_p,
    g472_n
  );


  or

  (
    g476_n,
    g453_n_spl_,
    g449_n_spl_
  );


  or

  (
    g477_n,
    g476_n_spl_,
    g457_n_spl_0
  );


  or

  (
    g478_n,
    g477_n,
    g461_p_spl_0
  );


  or

  (
    g479_n,
    g476_n_spl_,
    g457_p_spl_0
  );


  or

  (
    g480_n,
    g479_n,
    g461_n_spl_0
  );


  or

  (
    g481_n,
    g453_p_spl_0,
    g449_n_spl_
  );


  or

  (
    g482_n,
    g481_n,
    g457_n_spl_0
  );


  or

  (
    g483_n,
    g482_n,
    g461_n_spl_0
  );


  or

  (
    g484_n,
    g453_n_spl_,
    g449_p_spl_0
  );


  or

  (
    g485_n,
    g484_n,
    g457_n_spl_
  );


  or

  (
    g486_n,
    g485_n,
    g461_n_spl_
  );


  and

  (
    g487_p,
    g480_n,
    g478_n
  );


  and

  (
    g488_p,
    g487_p,
    g483_n
  );


  and

  (
    g489_p,
    g488_p,
    g486_n
  );


  and

  (
    g490_p,
    n1104_lo_p_spl_00,
    n1008_lo_p
  );


  or

  (
    g490_n,
    n1104_lo_n_spl_00,
    n1008_lo_n
  );


  and

  (
    g491_p,
    G627_o2_p_spl_0,
    G622_o2_p_spl_0
  );


  or

  (
    g491_n,
    G627_o2_n_spl_0,
    G622_o2_n_spl_0
  );


  and

  (
    g492_p,
    g491_n_spl_,
    G622_o2_p_spl_0
  );


  or

  (
    g492_n,
    g491_p_spl_,
    G622_o2_n_spl_0
  );


  and

  (
    g493_p,
    g491_n_spl_,
    G627_o2_p_spl_0
  );


  or

  (
    g493_n,
    g491_p_spl_,
    G627_o2_n_spl_0
  );


  and

  (
    g494_p,
    g493_n,
    g492_n
  );


  or

  (
    g494_n,
    g493_p,
    g492_p
  );


  and

  (
    g495_p,
    g494_n,
    g490_p
  );


  or

  (
    g496_n,
    g495_p_spl_,
    g490_n
  );


  or

  (
    g497_n,
    g495_p_spl_,
    g494_p
  );


  and

  (
    g498_p,
    g497_n,
    g496_n
  );


  and

  (
    g499_p,
    n1104_lo_p_spl_00,
    n1020_lo_p
  );


  or

  (
    g499_n,
    n1104_lo_n_spl_00,
    n1020_lo_n
  );


  and

  (
    g500_p,
    G637_o2_p_spl_0,
    G632_o2_p_spl_0
  );


  or

  (
    g500_n,
    G637_o2_n_spl_0,
    G632_o2_n_spl_0
  );


  and

  (
    g501_p,
    g500_n_spl_,
    G632_o2_p_spl_0
  );


  or

  (
    g501_n,
    g500_p_spl_,
    G632_o2_n_spl_0
  );


  and

  (
    g502_p,
    g500_n_spl_,
    G637_o2_p_spl_0
  );


  or

  (
    g502_n,
    g500_p_spl_,
    G637_o2_n_spl_0
  );


  and

  (
    g503_p,
    g502_n,
    g501_n
  );


  or

  (
    g503_n,
    g502_p,
    g501_p
  );


  and

  (
    g504_p,
    g503_n,
    g499_p
  );


  or

  (
    g505_n,
    g504_p_spl_,
    g499_n
  );


  or

  (
    g506_n,
    g504_p_spl_,
    g503_p
  );


  and

  (
    g507_p,
    g506_n,
    g505_n
  );


  and

  (
    g508_p,
    n1104_lo_p_spl_01,
    n1032_lo_p
  );


  or

  (
    g508_n,
    n1104_lo_n_spl_01,
    n1032_lo_n
  );


  and

  (
    g509_p,
    G632_o2_p_spl_1,
    G622_o2_p_spl_1
  );


  or

  (
    g509_n,
    G632_o2_n_spl_1,
    G622_o2_n_spl_1
  );


  and

  (
    g510_p,
    g509_n_spl_,
    G622_o2_p_spl_1
  );


  or

  (
    g510_n,
    g509_p_spl_,
    G622_o2_n_spl_1
  );


  and

  (
    g511_p,
    g509_n_spl_,
    G632_o2_p_spl_1
  );


  or

  (
    g511_n,
    g509_p_spl_,
    G632_o2_n_spl_1
  );


  and

  (
    g512_p,
    g511_n,
    g510_n
  );


  or

  (
    g512_n,
    g511_p,
    g510_p
  );


  and

  (
    g513_p,
    g512_n,
    g508_p
  );


  or

  (
    g514_n,
    g513_p_spl_,
    g508_n
  );


  or

  (
    g515_n,
    g513_p_spl_,
    g512_p
  );


  and

  (
    g516_p,
    g515_n,
    g514_n
  );


  and

  (
    g517_p,
    n1104_lo_p_spl_01,
    n1044_lo_p
  );


  or

  (
    g517_n,
    n1104_lo_n_spl_01,
    n1044_lo_n
  );


  and

  (
    g518_p,
    G637_o2_p_spl_1,
    G627_o2_p_spl_1
  );


  or

  (
    g518_n,
    G637_o2_n_spl_1,
    G627_o2_n_spl_1
  );


  and

  (
    g519_p,
    g518_n_spl_,
    G627_o2_p_spl_1
  );


  or

  (
    g519_n,
    g518_p_spl_,
    G627_o2_n_spl_1
  );


  and

  (
    g520_p,
    g518_n_spl_,
    G637_o2_p_spl_1
  );


  or

  (
    g520_n,
    g518_p_spl_,
    G637_o2_n_spl_1
  );


  and

  (
    g521_p,
    g520_n,
    g519_n
  );


  or

  (
    g521_n,
    g520_p,
    g519_p
  );


  and

  (
    g522_p,
    g521_n,
    g517_p
  );


  or

  (
    g523_n,
    g522_p_spl_,
    g517_n
  );


  or

  (
    g524_n,
    g522_p_spl_,
    g521_p
  );


  and

  (
    g525_p,
    g524_n,
    g523_n
  );


  and

  (
    g526_p,
    n1104_lo_p_spl_10,
    n1056_lo_p
  );


  or

  (
    g526_n,
    n1104_lo_n_spl_10,
    n1056_lo_n
  );


  and

  (
    g527_p,
    G607_o2_p_spl_0,
    G602_o2_p_spl_0
  );


  or

  (
    g527_n,
    G607_o2_n_spl_0,
    G602_o2_n_spl_0
  );


  and

  (
    g528_p,
    g527_n_spl_,
    G602_o2_p_spl_0
  );


  or

  (
    g528_n,
    g527_p_spl_,
    G602_o2_n_spl_0
  );


  and

  (
    g529_p,
    g527_n_spl_,
    G607_o2_p_spl_0
  );


  or

  (
    g529_n,
    g527_p_spl_,
    G607_o2_n_spl_0
  );


  and

  (
    g530_p,
    g529_n,
    g528_n
  );


  or

  (
    g530_n,
    g529_p,
    g528_p
  );


  and

  (
    g531_p,
    g530_n,
    g526_p
  );


  or

  (
    g532_n,
    g531_p_spl_,
    g526_n
  );


  or

  (
    g533_n,
    g531_p_spl_,
    g530_p
  );


  and

  (
    g534_p,
    g533_n,
    g532_n
  );


  and

  (
    g535_p,
    n1104_lo_p_spl_10,
    n1068_lo_p
  );


  or

  (
    g535_n,
    n1104_lo_n_spl_10,
    n1068_lo_n
  );


  and

  (
    g536_p,
    G617_o2_p_spl_0,
    G612_o2_p_spl_0
  );


  or

  (
    g536_n,
    G617_o2_n_spl_0,
    G612_o2_n_spl_0
  );


  and

  (
    g537_p,
    g536_n_spl_,
    G612_o2_p_spl_0
  );


  or

  (
    g537_n,
    g536_p_spl_,
    G612_o2_n_spl_0
  );


  and

  (
    g538_p,
    g536_n_spl_,
    G617_o2_p_spl_0
  );


  or

  (
    g538_n,
    g536_p_spl_,
    G617_o2_n_spl_0
  );


  and

  (
    g539_p,
    g538_n,
    g537_n
  );


  or

  (
    g539_n,
    g538_p,
    g537_p
  );


  and

  (
    g540_p,
    g539_n,
    g535_p
  );


  or

  (
    g541_n,
    g540_p_spl_,
    g535_n
  );


  or

  (
    g542_n,
    g540_p_spl_,
    g539_p
  );


  and

  (
    g543_p,
    g542_n,
    g541_n
  );


  and

  (
    g544_p,
    n1104_lo_p_spl_11,
    n1080_lo_p
  );


  or

  (
    g544_n,
    n1104_lo_n_spl_11,
    n1080_lo_n
  );


  and

  (
    g545_p,
    G612_o2_p_spl_1,
    G602_o2_p_spl_1
  );


  or

  (
    g545_n,
    G612_o2_n_spl_1,
    G602_o2_n_spl_1
  );


  and

  (
    g546_p,
    g545_n_spl_,
    G602_o2_p_spl_1
  );


  or

  (
    g546_n,
    g545_p_spl_,
    G602_o2_n_spl_1
  );


  and

  (
    g547_p,
    g545_n_spl_,
    G612_o2_p_spl_1
  );


  or

  (
    g547_n,
    g545_p_spl_,
    G612_o2_n_spl_1
  );


  and

  (
    g548_p,
    g547_n,
    g546_n
  );


  or

  (
    g548_n,
    g547_p,
    g546_p
  );


  and

  (
    g549_p,
    g548_n,
    g544_p
  );


  or

  (
    g550_n,
    g549_p_spl_,
    g544_n
  );


  or

  (
    g551_n,
    g549_p_spl_,
    g548_p
  );


  and

  (
    g552_p,
    g551_n,
    g550_n
  );


  and

  (
    g553_p,
    n1104_lo_p_spl_11,
    n1092_lo_p
  );


  or

  (
    g553_n,
    n1104_lo_n_spl_11,
    n1092_lo_n
  );


  and

  (
    g554_p,
    G617_o2_p_spl_1,
    G607_o2_p_spl_1
  );


  or

  (
    g554_n,
    G617_o2_n_spl_1,
    G607_o2_n_spl_1
  );


  and

  (
    g555_p,
    g554_n_spl_,
    G607_o2_p_spl_1
  );


  or

  (
    g555_n,
    g554_p_spl_,
    G607_o2_n_spl_1
  );


  and

  (
    g556_p,
    g554_n_spl_,
    G617_o2_p_spl_1
  );


  or

  (
    g556_n,
    g554_p_spl_,
    G617_o2_n_spl_1
  );


  and

  (
    g557_p,
    g556_n,
    g555_n
  );


  or

  (
    g557_n,
    g556_p,
    g555_p
  );


  and

  (
    g558_p,
    g557_n,
    g553_p
  );


  or

  (
    g559_n,
    g558_p_spl_,
    g553_n
  );


  or

  (
    g560_n,
    g558_p_spl_,
    g557_p
  );


  and

  (
    g561_p,
    g560_n,
    g559_n
  );


  and

  (
    g562_p,
    n2155_o2_p_spl_,
    n2151_o2_p_spl_
  );


  or

  (
    g562_n,
    n2155_o2_n_spl_0,
    n2151_o2_n_spl_0
  );


  and

  (
    g563_p,
    g562_n_spl_,
    n2151_o2_p_spl_
  );


  or

  (
    g563_n,
    g562_p_spl_,
    n2151_o2_n_spl_0
  );


  and

  (
    g564_p,
    g562_n_spl_,
    n2155_o2_p_spl_
  );


  or

  (
    g564_n,
    g562_p_spl_,
    n2155_o2_n_spl_0
  );


  and

  (
    g565_p,
    g564_n,
    g563_n
  );


  or

  (
    g565_n,
    g564_p,
    g563_p
  );


  and

  (
    g566_p,
    n2163_o2_p_spl_,
    n2159_o2_p_spl_
  );


  or

  (
    g566_n,
    n2163_o2_n_spl_0,
    n2159_o2_n_spl_0
  );


  and

  (
    g567_p,
    g566_n_spl_,
    n2159_o2_p_spl_
  );


  or

  (
    g567_n,
    g566_p_spl_,
    n2159_o2_n_spl_0
  );


  and

  (
    g568_p,
    g566_n_spl_,
    n2163_o2_p_spl_
  );


  or

  (
    g568_n,
    g566_p_spl_,
    n2163_o2_n_spl_0
  );


  and

  (
    g569_p,
    g568_n,
    g567_n
  );


  or

  (
    g569_n,
    g568_p,
    g567_p
  );


  and

  (
    g570_p,
    g569_n,
    g565_n
  );


  or

  (
    g571_n,
    g570_p_spl_,
    g565_p
  );


  or

  (
    g572_n,
    g570_p_spl_,
    g569_p
  );


  and

  (
    g573_p,
    g572_n,
    g571_n
  );


  and

  (
    g574_p,
    n2156_o2_p_spl_,
    n2152_o2_p_spl_
  );


  or

  (
    g574_n,
    n2156_o2_n_spl_0,
    n2152_o2_n_spl_0
  );


  and

  (
    g575_p,
    g574_n_spl_,
    n2152_o2_p_spl_
  );


  or

  (
    g575_n,
    g574_p_spl_,
    n2152_o2_n_spl_0
  );


  and

  (
    g576_p,
    g574_n_spl_,
    n2156_o2_p_spl_
  );


  or

  (
    g576_n,
    g574_p_spl_,
    n2156_o2_n_spl_0
  );


  and

  (
    g577_p,
    g576_n,
    g575_n
  );


  or

  (
    g577_n,
    g576_p,
    g575_p
  );


  and

  (
    g578_p,
    n2164_o2_p_spl_,
    n2160_o2_p_spl_
  );


  or

  (
    g578_n,
    n2164_o2_n_spl_0,
    n2160_o2_n_spl_0
  );


  and

  (
    g579_p,
    g578_n_spl_,
    n2160_o2_p_spl_
  );


  or

  (
    g579_n,
    g578_p_spl_,
    n2160_o2_n_spl_0
  );


  and

  (
    g580_p,
    g578_n_spl_,
    n2164_o2_p_spl_
  );


  or

  (
    g580_n,
    g578_p_spl_,
    n2164_o2_n_spl_0
  );


  and

  (
    g581_p,
    g580_n,
    g579_n
  );


  or

  (
    g581_n,
    g580_p,
    g579_p
  );


  and

  (
    g582_p,
    g581_n,
    g577_n
  );


  or

  (
    g583_n,
    g582_p_spl_,
    g577_p
  );


  or

  (
    g584_n,
    g582_p_spl_,
    g581_p
  );


  and

  (
    g585_p,
    g584_n,
    g583_n
  );


  and

  (
    g586_p,
    n2157_o2_p_spl_,
    n2153_o2_p_spl_
  );


  or

  (
    g586_n,
    n2157_o2_n_spl_0,
    n2153_o2_n_spl_0
  );


  and

  (
    g587_p,
    g586_n_spl_,
    n2153_o2_p_spl_
  );


  or

  (
    g587_n,
    g586_p_spl_,
    n2153_o2_n_spl_0
  );


  and

  (
    g588_p,
    g586_n_spl_,
    n2157_o2_p_spl_
  );


  or

  (
    g588_n,
    g586_p_spl_,
    n2157_o2_n_spl_0
  );


  and

  (
    g589_p,
    g588_n,
    g587_n
  );


  or

  (
    g589_n,
    g588_p,
    g587_p
  );


  and

  (
    g590_p,
    n2165_o2_p_spl_,
    n2161_o2_p_spl_
  );


  or

  (
    g590_n,
    n2165_o2_n_spl_0,
    n2161_o2_n_spl_0
  );


  and

  (
    g591_p,
    g590_n_spl_,
    n2161_o2_p_spl_
  );


  or

  (
    g591_n,
    g590_p_spl_,
    n2161_o2_n_spl_0
  );


  and

  (
    g592_p,
    g590_n_spl_,
    n2165_o2_p_spl_
  );


  or

  (
    g592_n,
    g590_p_spl_,
    n2165_o2_n_spl_0
  );


  and

  (
    g593_p,
    g592_n,
    g591_n
  );


  or

  (
    g593_n,
    g592_p,
    g591_p
  );


  and

  (
    g594_p,
    g593_n,
    g589_n
  );


  or

  (
    g595_n,
    g594_p_spl_,
    g589_p
  );


  or

  (
    g596_n,
    g594_p_spl_,
    g593_p
  );


  and

  (
    g597_p,
    g596_n,
    g595_n
  );


  and

  (
    g598_p,
    n2158_o2_p_spl_,
    n2154_o2_p_spl_
  );


  or

  (
    g598_n,
    n2158_o2_n_spl_0,
    n2154_o2_n_spl_0
  );


  and

  (
    g599_p,
    g598_n_spl_,
    n2154_o2_p_spl_
  );


  or

  (
    g599_n,
    g598_p_spl_,
    n2154_o2_n_spl_0
  );


  and

  (
    g600_p,
    g598_n_spl_,
    n2158_o2_p_spl_
  );


  or

  (
    g600_n,
    g598_p_spl_,
    n2158_o2_n_spl_0
  );


  and

  (
    g601_p,
    g600_n,
    g599_n
  );


  or

  (
    g601_n,
    g600_p,
    g599_p
  );


  and

  (
    g602_p,
    n2166_o2_p_spl_,
    n2162_o2_p_spl_
  );


  or

  (
    g602_n,
    n2166_o2_n_spl_0,
    n2162_o2_n_spl_0
  );


  and

  (
    g603_p,
    g602_n_spl_,
    n2162_o2_p_spl_
  );


  or

  (
    g603_n,
    g602_p_spl_,
    n2162_o2_n_spl_0
  );


  and

  (
    g604_p,
    g602_n_spl_,
    n2166_o2_p_spl_
  );


  or

  (
    g604_n,
    g602_p_spl_,
    n2166_o2_n_spl_0
  );


  and

  (
    g605_p,
    g604_n,
    g603_n
  );


  or

  (
    g605_n,
    g604_p,
    g603_p
  );


  and

  (
    g606_p,
    g605_n,
    g601_n
  );


  or

  (
    g607_n,
    g606_p_spl_,
    g601_p
  );


  or

  (
    g608_n,
    g606_p_spl_,
    g605_p
  );


  and

  (
    g609_p,
    g608_n,
    g607_n
  );


  and

  (
    g610_p,
    n2171_o2_p_spl_,
    n2167_o2_p_spl_
  );


  or

  (
    g610_n,
    n2171_o2_n_spl_0,
    n2167_o2_n_spl_0
  );


  and

  (
    g611_p,
    g610_n_spl_,
    n2167_o2_p_spl_
  );


  or

  (
    g611_n,
    g610_p_spl_,
    n2167_o2_n_spl_0
  );


  and

  (
    g612_p,
    g610_n_spl_,
    n2171_o2_p_spl_
  );


  or

  (
    g612_n,
    g610_p_spl_,
    n2171_o2_n_spl_0
  );


  and

  (
    g613_p,
    g612_n,
    g611_n
  );


  or

  (
    g613_n,
    g612_p,
    g611_p
  );


  and

  (
    g614_p,
    n2179_o2_p_spl_,
    n2175_o2_p_spl_
  );


  or

  (
    g614_n,
    n2179_o2_n_spl_0,
    n2175_o2_n_spl_0
  );


  and

  (
    g615_p,
    g614_n_spl_,
    n2175_o2_p_spl_
  );


  or

  (
    g615_n,
    g614_p_spl_,
    n2175_o2_n_spl_0
  );


  and

  (
    g616_p,
    g614_n_spl_,
    n2179_o2_p_spl_
  );


  or

  (
    g616_n,
    g614_p_spl_,
    n2179_o2_n_spl_0
  );


  and

  (
    g617_p,
    g616_n,
    g615_n
  );


  or

  (
    g617_n,
    g616_p,
    g615_p
  );


  and

  (
    g618_p,
    g617_n,
    g613_n
  );


  or

  (
    g619_n,
    g618_p_spl_,
    g613_p
  );


  or

  (
    g620_n,
    g618_p_spl_,
    g617_p
  );


  and

  (
    g621_p,
    g620_n,
    g619_n
  );


  and

  (
    g622_p,
    n2172_o2_p_spl_,
    n2168_o2_p_spl_
  );


  or

  (
    g622_n,
    n2172_o2_n_spl_0,
    n2168_o2_n_spl_0
  );


  and

  (
    g623_p,
    g622_n_spl_,
    n2168_o2_p_spl_
  );


  or

  (
    g623_n,
    g622_p_spl_,
    n2168_o2_n_spl_0
  );


  and

  (
    g624_p,
    g622_n_spl_,
    n2172_o2_p_spl_
  );


  or

  (
    g624_n,
    g622_p_spl_,
    n2172_o2_n_spl_0
  );


  and

  (
    g625_p,
    g624_n,
    g623_n
  );


  or

  (
    g625_n,
    g624_p,
    g623_p
  );


  and

  (
    g626_p,
    n2180_o2_p_spl_,
    n2176_o2_p_spl_
  );


  or

  (
    g626_n,
    n2180_o2_n_spl_0,
    n2176_o2_n_spl_0
  );


  and

  (
    g627_p,
    g626_n_spl_,
    n2176_o2_p_spl_
  );


  or

  (
    g627_n,
    g626_p_spl_,
    n2176_o2_n_spl_0
  );


  and

  (
    g628_p,
    g626_n_spl_,
    n2180_o2_p_spl_
  );


  or

  (
    g628_n,
    g626_p_spl_,
    n2180_o2_n_spl_0
  );


  and

  (
    g629_p,
    g628_n,
    g627_n
  );


  or

  (
    g629_n,
    g628_p,
    g627_p
  );


  and

  (
    g630_p,
    g629_n,
    g625_n
  );


  or

  (
    g631_n,
    g630_p_spl_,
    g625_p
  );


  or

  (
    g632_n,
    g630_p_spl_,
    g629_p
  );


  and

  (
    g633_p,
    g632_n,
    g631_n
  );


  and

  (
    g634_p,
    n2173_o2_p_spl_,
    n2169_o2_p_spl_
  );


  or

  (
    g634_n,
    n2173_o2_n_spl_0,
    n2169_o2_n_spl_0
  );


  and

  (
    g635_p,
    g634_n_spl_,
    n2169_o2_p_spl_
  );


  or

  (
    g635_n,
    g634_p_spl_,
    n2169_o2_n_spl_0
  );


  and

  (
    g636_p,
    g634_n_spl_,
    n2173_o2_p_spl_
  );


  or

  (
    g636_n,
    g634_p_spl_,
    n2173_o2_n_spl_0
  );


  and

  (
    g637_p,
    g636_n,
    g635_n
  );


  or

  (
    g637_n,
    g636_p,
    g635_p
  );


  and

  (
    g638_p,
    n2181_o2_p_spl_,
    n2177_o2_p_spl_
  );


  or

  (
    g638_n,
    n2181_o2_n_spl_0,
    n2177_o2_n_spl_0
  );


  and

  (
    g639_p,
    g638_n_spl_,
    n2177_o2_p_spl_
  );


  or

  (
    g639_n,
    g638_p_spl_,
    n2177_o2_n_spl_0
  );


  and

  (
    g640_p,
    g638_n_spl_,
    n2181_o2_p_spl_
  );


  or

  (
    g640_n,
    g638_p_spl_,
    n2181_o2_n_spl_0
  );


  and

  (
    g641_p,
    g640_n,
    g639_n
  );


  or

  (
    g641_n,
    g640_p,
    g639_p
  );


  and

  (
    g642_p,
    g641_n,
    g637_n
  );


  or

  (
    g643_n,
    g642_p_spl_,
    g637_p
  );


  or

  (
    g644_n,
    g642_p_spl_,
    g641_p
  );


  and

  (
    g645_p,
    g644_n,
    g643_n
  );


  and

  (
    g646_p,
    n2174_o2_p_spl_,
    n2170_o2_p_spl_
  );


  or

  (
    g646_n,
    n2174_o2_n_spl_0,
    n2170_o2_n_spl_0
  );


  and

  (
    g647_p,
    g646_n_spl_,
    n2170_o2_p_spl_
  );


  or

  (
    g647_n,
    g646_p_spl_,
    n2170_o2_n_spl_0
  );


  and

  (
    g648_p,
    g646_n_spl_,
    n2174_o2_p_spl_
  );


  or

  (
    g648_n,
    g646_p_spl_,
    n2174_o2_n_spl_0
  );


  and

  (
    g649_p,
    g648_n,
    g647_n
  );


  or

  (
    g649_n,
    g648_p,
    g647_p
  );


  and

  (
    g650_p,
    n2182_o2_p_spl_,
    n2178_o2_p_spl_
  );


  or

  (
    g650_n,
    n2182_o2_n_spl_0,
    n2178_o2_n_spl_0
  );


  and

  (
    g651_p,
    g650_n_spl_,
    n2178_o2_p_spl_
  );


  or

  (
    g651_n,
    g650_p_spl_,
    n2178_o2_n_spl_0
  );


  and

  (
    g652_p,
    g650_n_spl_,
    n2182_o2_p_spl_
  );


  or

  (
    g652_n,
    g650_p_spl_,
    n2182_o2_n_spl_0
  );


  and

  (
    g653_p,
    g652_n,
    g651_n
  );


  or

  (
    g653_n,
    g652_p,
    g651_p
  );


  and

  (
    g654_p,
    g653_n,
    g649_n
  );


  or

  (
    g655_n,
    g654_p_spl_,
    g649_p
  );


  or

  (
    g656_n,
    g654_p_spl_,
    g653_p
  );


  and

  (
    g657_p,
    g656_n,
    g655_n
  );


  and

  (
    g658_p,
    n639_lo_buf_o2_p_spl_,
    n627_lo_buf_o2_p_spl_
  );


  or

  (
    g658_n,
    n639_lo_buf_o2_n_spl_0,
    n627_lo_buf_o2_n_spl_0
  );


  and

  (
    g659_p,
    g658_n_spl_,
    n627_lo_buf_o2_p_spl_
  );


  or

  (
    g659_n,
    g658_p_spl_,
    n627_lo_buf_o2_n_spl_0
  );


  and

  (
    g660_p,
    g658_n_spl_,
    n639_lo_buf_o2_p_spl_
  );


  or

  (
    g660_n,
    g658_p_spl_,
    n639_lo_buf_o2_n_spl_0
  );


  and

  (
    g661_p,
    g660_n,
    g659_n
  );


  or

  (
    g661_n,
    g660_p,
    g659_p
  );


  and

  (
    g662_p,
    n663_lo_buf_o2_p_spl_,
    n651_lo_buf_o2_p_spl_
  );


  or

  (
    g662_n,
    n663_lo_buf_o2_n_spl_0,
    n651_lo_buf_o2_n_spl_0
  );


  and

  (
    g663_p,
    g662_n_spl_,
    n651_lo_buf_o2_p_spl_
  );


  or

  (
    g663_n,
    g662_p_spl_,
    n651_lo_buf_o2_n_spl_0
  );


  and

  (
    g664_p,
    g662_n_spl_,
    n663_lo_buf_o2_p_spl_
  );


  or

  (
    g664_n,
    g662_p_spl_,
    n663_lo_buf_o2_n_spl_0
  );


  and

  (
    g665_p,
    g664_n,
    g663_n
  );


  or

  (
    g665_n,
    g664_p,
    g663_p
  );


  and

  (
    g666_p,
    g665_n,
    g661_n
  );


  or

  (
    g667_n,
    g666_p_spl_,
    g661_p
  );


  or

  (
    g668_n,
    g666_p_spl_,
    g665_p
  );


  and

  (
    g669_p,
    g668_n,
    g667_n
  );


  and

  (
    g670_p,
    n687_lo_buf_o2_p_spl_,
    n675_lo_buf_o2_p_spl_
  );


  or

  (
    g670_n,
    n687_lo_buf_o2_n_spl_0,
    n675_lo_buf_o2_n_spl_0
  );


  and

  (
    g671_p,
    g670_n_spl_,
    n675_lo_buf_o2_p_spl_
  );


  or

  (
    g671_n,
    g670_p_spl_,
    n675_lo_buf_o2_n_spl_0
  );


  and

  (
    g672_p,
    g670_n_spl_,
    n687_lo_buf_o2_p_spl_
  );


  or

  (
    g672_n,
    g670_p_spl_,
    n687_lo_buf_o2_n_spl_0
  );


  and

  (
    g673_p,
    g672_n,
    g671_n
  );


  or

  (
    g673_n,
    g672_p,
    g671_p
  );


  and

  (
    g674_p,
    n711_lo_buf_o2_p_spl_,
    n699_lo_buf_o2_p_spl_
  );


  or

  (
    g674_n,
    n711_lo_buf_o2_n_spl_0,
    n699_lo_buf_o2_n_spl_0
  );


  and

  (
    g675_p,
    g674_n_spl_,
    n699_lo_buf_o2_p_spl_
  );


  or

  (
    g675_n,
    g674_p_spl_,
    n699_lo_buf_o2_n_spl_0
  );


  and

  (
    g676_p,
    g674_n_spl_,
    n711_lo_buf_o2_p_spl_
  );


  or

  (
    g676_n,
    g674_p_spl_,
    n711_lo_buf_o2_n_spl_0
  );


  and

  (
    g677_p,
    g676_n,
    g675_n
  );


  or

  (
    g677_n,
    g676_p,
    g675_p
  );


  and

  (
    g678_p,
    g677_n,
    g673_n
  );


  or

  (
    g679_n,
    g678_p_spl_,
    g673_p
  );


  or

  (
    g680_n,
    g678_p_spl_,
    g677_p
  );


  and

  (
    g681_p,
    g680_n,
    g679_n
  );


  and

  (
    g682_p,
    n735_lo_buf_o2_p_spl_,
    n723_lo_buf_o2_p_spl_
  );


  or

  (
    g682_n,
    n735_lo_buf_o2_n_spl_0,
    n723_lo_buf_o2_n_spl_0
  );


  and

  (
    g683_p,
    g682_n_spl_,
    n723_lo_buf_o2_p_spl_
  );


  or

  (
    g683_n,
    g682_p_spl_,
    n723_lo_buf_o2_n_spl_0
  );


  and

  (
    g684_p,
    g682_n_spl_,
    n735_lo_buf_o2_p_spl_
  );


  or

  (
    g684_n,
    g682_p_spl_,
    n735_lo_buf_o2_n_spl_0
  );


  and

  (
    g685_p,
    g684_n,
    g683_n
  );


  or

  (
    g685_n,
    g684_p,
    g683_p
  );


  and

  (
    g686_p,
    n759_lo_buf_o2_p_spl_,
    n747_lo_buf_o2_p_spl_
  );


  or

  (
    g686_n,
    n759_lo_buf_o2_n_spl_0,
    n747_lo_buf_o2_n_spl_0
  );


  and

  (
    g687_p,
    g686_n_spl_,
    n747_lo_buf_o2_p_spl_
  );


  or

  (
    g687_n,
    g686_p_spl_,
    n747_lo_buf_o2_n_spl_0
  );


  and

  (
    g688_p,
    g686_n_spl_,
    n759_lo_buf_o2_p_spl_
  );


  or

  (
    g688_n,
    g686_p_spl_,
    n759_lo_buf_o2_n_spl_0
  );


  and

  (
    g689_p,
    g688_n,
    g687_n
  );


  or

  (
    g689_n,
    g688_p,
    g687_p
  );


  and

  (
    g690_p,
    g689_n,
    g685_n
  );


  or

  (
    g691_n,
    g690_p_spl_,
    g685_p
  );


  or

  (
    g692_n,
    g690_p_spl_,
    g689_p
  );


  and

  (
    g693_p,
    g692_n,
    g691_n
  );


  and

  (
    g694_p,
    n783_lo_buf_o2_p_spl_,
    n771_lo_buf_o2_p_spl_
  );


  or

  (
    g694_n,
    n783_lo_buf_o2_n_spl_0,
    n771_lo_buf_o2_n_spl_0
  );


  and

  (
    g695_p,
    g694_n_spl_,
    n771_lo_buf_o2_p_spl_
  );


  or

  (
    g695_n,
    g694_p_spl_,
    n771_lo_buf_o2_n_spl_0
  );


  and

  (
    g696_p,
    g694_n_spl_,
    n783_lo_buf_o2_p_spl_
  );


  or

  (
    g696_n,
    g694_p_spl_,
    n783_lo_buf_o2_n_spl_0
  );


  and

  (
    g697_p,
    g696_n,
    g695_n
  );


  or

  (
    g697_n,
    g696_p,
    g695_p
  );


  and

  (
    g698_p,
    n807_lo_buf_o2_p_spl_,
    n795_lo_buf_o2_p_spl_
  );


  or

  (
    g698_n,
    n807_lo_buf_o2_n_spl_0,
    n795_lo_buf_o2_n_spl_0
  );


  and

  (
    g699_p,
    g698_n_spl_,
    n795_lo_buf_o2_p_spl_
  );


  or

  (
    g699_n,
    g698_p_spl_,
    n795_lo_buf_o2_n_spl_0
  );


  and

  (
    g700_p,
    g698_n_spl_,
    n807_lo_buf_o2_p_spl_
  );


  or

  (
    g700_n,
    g698_p_spl_,
    n807_lo_buf_o2_n_spl_0
  );


  and

  (
    g701_p,
    g700_n,
    g699_n
  );


  or

  (
    g701_n,
    g700_p,
    g699_p
  );


  and

  (
    g702_p,
    g701_n,
    g697_n
  );


  or

  (
    g703_n,
    g702_p_spl_,
    g697_p
  );


  or

  (
    g704_n,
    g702_p_spl_,
    g701_p
  );


  and

  (
    g705_p,
    g704_n,
    g703_n
  );


  and

  (
    g706_p,
    n831_lo_buf_o2_p_spl_,
    n819_lo_buf_o2_p_spl_
  );


  or

  (
    g706_n,
    n831_lo_buf_o2_n_spl_0,
    n819_lo_buf_o2_n_spl_0
  );


  and

  (
    g707_p,
    g706_n_spl_,
    n819_lo_buf_o2_p_spl_
  );


  or

  (
    g707_n,
    g706_p_spl_,
    n819_lo_buf_o2_n_spl_0
  );


  and

  (
    g708_p,
    g706_n_spl_,
    n831_lo_buf_o2_p_spl_
  );


  or

  (
    g708_n,
    g706_p_spl_,
    n831_lo_buf_o2_n_spl_0
  );


  and

  (
    g709_p,
    g708_n,
    g707_n
  );


  or

  (
    g709_n,
    g708_p,
    g707_p
  );


  and

  (
    g710_p,
    n855_lo_buf_o2_p_spl_,
    n843_lo_buf_o2_p_spl_
  );


  or

  (
    g710_n,
    n855_lo_buf_o2_n_spl_0,
    n843_lo_buf_o2_n_spl_0
  );


  and

  (
    g711_p,
    g710_n_spl_,
    n843_lo_buf_o2_p_spl_
  );


  or

  (
    g711_n,
    g710_p_spl_,
    n843_lo_buf_o2_n_spl_0
  );


  and

  (
    g712_p,
    g710_n_spl_,
    n855_lo_buf_o2_p_spl_
  );


  or

  (
    g712_n,
    g710_p_spl_,
    n855_lo_buf_o2_n_spl_0
  );


  and

  (
    g713_p,
    g712_n,
    g711_n
  );


  or

  (
    g713_n,
    g712_p,
    g711_p
  );


  and

  (
    g714_p,
    g713_n,
    g709_n
  );


  or

  (
    g715_n,
    g714_p_spl_,
    g709_p
  );


  or

  (
    g716_n,
    g714_p_spl_,
    g713_p
  );


  and

  (
    g717_p,
    g716_n,
    g715_n
  );


  and

  (
    g718_p,
    n879_lo_buf_o2_p_spl_,
    n867_lo_buf_o2_p_spl_
  );


  or

  (
    g718_n,
    n879_lo_buf_o2_n_spl_0,
    n867_lo_buf_o2_n_spl_0
  );


  and

  (
    g719_p,
    g718_n_spl_,
    n867_lo_buf_o2_p_spl_
  );


  or

  (
    g719_n,
    g718_p_spl_,
    n867_lo_buf_o2_n_spl_0
  );


  and

  (
    g720_p,
    g718_n_spl_,
    n879_lo_buf_o2_p_spl_
  );


  or

  (
    g720_n,
    g718_p_spl_,
    n879_lo_buf_o2_n_spl_0
  );


  and

  (
    g721_p,
    g720_n,
    g719_n
  );


  or

  (
    g721_n,
    g720_p,
    g719_p
  );


  and

  (
    g722_p,
    n903_lo_buf_o2_p_spl_,
    n891_lo_buf_o2_p_spl_
  );


  or

  (
    g722_n,
    n903_lo_buf_o2_n_spl_0,
    n891_lo_buf_o2_n_spl_0
  );


  and

  (
    g723_p,
    g722_n_spl_,
    n891_lo_buf_o2_p_spl_
  );


  or

  (
    g723_n,
    g722_p_spl_,
    n891_lo_buf_o2_n_spl_0
  );


  and

  (
    g724_p,
    g722_n_spl_,
    n903_lo_buf_o2_p_spl_
  );


  or

  (
    g724_n,
    g722_p_spl_,
    n903_lo_buf_o2_n_spl_0
  );


  and

  (
    g725_p,
    g724_n,
    g723_n
  );


  or

  (
    g725_n,
    g724_p,
    g723_p
  );


  and

  (
    g726_p,
    g725_n,
    g721_n
  );


  or

  (
    g727_n,
    g726_p_spl_,
    g721_p
  );


  or

  (
    g728_n,
    g726_p_spl_,
    g725_p
  );


  and

  (
    g729_p,
    g728_n,
    g727_n
  );


  and

  (
    g730_p,
    n927_lo_buf_o2_p_spl_,
    n915_lo_buf_o2_p_spl_
  );


  or

  (
    g730_n,
    n927_lo_buf_o2_n_spl_0,
    n915_lo_buf_o2_n_spl_0
  );


  and

  (
    g731_p,
    g730_n_spl_,
    n915_lo_buf_o2_p_spl_
  );


  or

  (
    g731_n,
    g730_p_spl_,
    n915_lo_buf_o2_n_spl_0
  );


  and

  (
    g732_p,
    g730_n_spl_,
    n927_lo_buf_o2_p_spl_
  );


  or

  (
    g732_n,
    g730_p_spl_,
    n927_lo_buf_o2_n_spl_0
  );


  and

  (
    g733_p,
    g732_n,
    g731_n
  );


  or

  (
    g733_n,
    g732_p,
    g731_p
  );


  and

  (
    g734_p,
    n951_lo_buf_o2_p_spl_,
    n939_lo_buf_o2_p_spl_
  );


  or

  (
    g734_n,
    n951_lo_buf_o2_n_spl_0,
    n939_lo_buf_o2_n_spl_0
  );


  and

  (
    g735_p,
    g734_n_spl_,
    n939_lo_buf_o2_p_spl_
  );


  or

  (
    g735_n,
    g734_p_spl_,
    n939_lo_buf_o2_n_spl_0
  );


  and

  (
    g736_p,
    g734_n_spl_,
    n951_lo_buf_o2_p_spl_
  );


  or

  (
    g736_n,
    g734_p_spl_,
    n951_lo_buf_o2_n_spl_0
  );


  and

  (
    g737_p,
    g736_n,
    g735_n
  );


  or

  (
    g737_n,
    g736_p,
    g735_p
  );


  and

  (
    g738_p,
    g737_n,
    g733_n
  );


  or

  (
    g739_n,
    g738_p_spl_,
    g733_p
  );


  or

  (
    g740_n,
    g738_p_spl_,
    g737_p
  );


  and

  (
    g741_p,
    g740_n,
    g739_n
  );


  and

  (
    g742_p,
    n975_lo_buf_o2_p_spl_,
    n963_lo_buf_o2_p_spl_
  );


  or

  (
    g742_n,
    n975_lo_buf_o2_n_spl_0,
    n963_lo_buf_o2_n_spl_0
  );


  and

  (
    g743_p,
    g742_n_spl_,
    n963_lo_buf_o2_p_spl_
  );


  or

  (
    g743_n,
    g742_p_spl_,
    n963_lo_buf_o2_n_spl_0
  );


  and

  (
    g744_p,
    g742_n_spl_,
    n975_lo_buf_o2_p_spl_
  );


  or

  (
    g744_n,
    g742_p_spl_,
    n975_lo_buf_o2_n_spl_0
  );


  and

  (
    g745_p,
    g744_n,
    g743_n
  );


  or

  (
    g745_n,
    g744_p,
    g743_p
  );


  and

  (
    g746_p,
    n999_lo_buf_o2_p_spl_,
    n987_lo_buf_o2_p_spl_
  );


  or

  (
    g746_n,
    n999_lo_buf_o2_n_spl_0,
    n987_lo_buf_o2_n_spl_0
  );


  and

  (
    g747_p,
    g746_n_spl_,
    n987_lo_buf_o2_p_spl_
  );


  or

  (
    g747_n,
    g746_p_spl_,
    n987_lo_buf_o2_n_spl_0
  );


  and

  (
    g748_p,
    g746_n_spl_,
    n999_lo_buf_o2_p_spl_
  );


  or

  (
    g748_n,
    g746_p_spl_,
    n999_lo_buf_o2_n_spl_0
  );


  and

  (
    g749_p,
    g748_n,
    g747_n
  );


  or

  (
    g749_n,
    g748_p,
    g747_p
  );


  and

  (
    g750_p,
    g749_n,
    g745_n
  );


  or

  (
    g751_n,
    g750_p_spl_,
    g745_p
  );


  or

  (
    g752_n,
    g750_p_spl_,
    g749_p
  );


  and

  (
    g753_p,
    g752_n,
    g751_n
  );


  not

  (
    G1324,
    g246_n
  );


  not

  (
    G1325,
    g251_n
  );


  not

  (
    G1326,
    g256_n
  );


  not

  (
    G1327,
    g261_n
  );


  not

  (
    G1328,
    g270_n
  );


  not

  (
    G1329,
    g275_n
  );


  not

  (
    G1330,
    g280_n
  );


  not

  (
    G1331,
    g285_n
  );


  not

  (
    G1332,
    g294_n
  );


  not

  (
    G1333,
    g299_n
  );


  not

  (
    G1334,
    g304_n
  );


  not

  (
    G1335,
    g309_n
  );


  not

  (
    G1336,
    g318_n
  );


  not

  (
    G1337,
    g323_n
  );


  not

  (
    G1338,
    g328_n
  );


  not

  (
    G1339,
    g333_n
  );


  not

  (
    G1340,
    g342_n
  );


  not

  (
    G1341,
    g347_n
  );


  not

  (
    G1342,
    g352_n
  );


  not

  (
    G1343,
    g357_n
  );


  not

  (
    G1344,
    g366_n
  );


  not

  (
    G1345,
    g371_n
  );


  not

  (
    G1346,
    g376_n
  );


  not

  (
    G1347,
    g381_n
  );


  not

  (
    G1348,
    g390_n
  );


  not

  (
    G1349,
    g395_n
  );


  not

  (
    G1350,
    g400_n
  );


  not

  (
    G1351,
    g405_n
  );


  not

  (
    G1352,
    g414_n
  );


  not

  (
    G1353,
    g419_n
  );


  not

  (
    G1354,
    g424_n
  );


  not

  (
    G1355,
    g429_n
  );


  not

  (
    n630_li,
    n1837_o2_n
  );


  not

  (
    n642_li,
    n1838_o2_n
  );


  not

  (
    n654_li,
    n1839_o2_n
  );


  not

  (
    n666_li,
    n1840_o2_n
  );


  not

  (
    n678_li,
    n1841_o2_n
  );


  not

  (
    n690_li,
    n1842_o2_n
  );


  not

  (
    n702_li,
    n1843_o2_n
  );


  not

  (
    n714_li,
    n1844_o2_n
  );


  not

  (
    n726_li,
    n1845_o2_n
  );


  not

  (
    n738_li,
    n1846_o2_n
  );


  not

  (
    n750_li,
    n1847_o2_n
  );


  not

  (
    n762_li,
    n1848_o2_n
  );


  not

  (
    n774_li,
    n1849_o2_n
  );


  not

  (
    n786_li,
    n1850_o2_n
  );


  not

  (
    n798_li,
    n1851_o2_n
  );


  not

  (
    n810_li,
    n1852_o2_n
  );


  not

  (
    n822_li,
    n1853_o2_n
  );


  not

  (
    n834_li,
    n1854_o2_n
  );


  not

  (
    n846_li,
    n1855_o2_n
  );


  not

  (
    n858_li,
    n1856_o2_n
  );


  not

  (
    n870_li,
    n1857_o2_n
  );


  not

  (
    n882_li,
    n1858_o2_n
  );


  not

  (
    n894_li,
    n1859_o2_n
  );


  not

  (
    n906_li,
    n1860_o2_n
  );


  not

  (
    n918_li,
    n1861_o2_n
  );


  not

  (
    n930_li,
    n1862_o2_n
  );


  not

  (
    n942_li,
    n1863_o2_n
  );


  not

  (
    n954_li,
    n1864_o2_n
  );


  not

  (
    n966_li,
    n1865_o2_n
  );


  not

  (
    n978_li,
    n1866_o2_n
  );


  not

  (
    n990_li,
    n1867_o2_n
  );


  not

  (
    n1002_li,
    n1868_o2_n
  );


  not

  (
    n1005_li,
    G33_n
  );


  not

  (
    n1008_li,
    n1005_lo_n
  );


  not

  (
    n1017_li,
    G34_n
  );


  not

  (
    n1020_li,
    n1017_lo_n
  );


  not

  (
    n1029_li,
    G35_n
  );


  not

  (
    n1032_li,
    n1029_lo_n
  );


  not

  (
    n1041_li,
    G36_n
  );


  not

  (
    n1044_li,
    n1041_lo_n
  );


  not

  (
    n1053_li,
    G37_n
  );


  not

  (
    n1056_li,
    n1053_lo_n
  );


  not

  (
    n1065_li,
    G38_n
  );


  not

  (
    n1068_li,
    n1065_lo_n
  );


  not

  (
    n1077_li,
    G39_n
  );


  not

  (
    n1080_li,
    n1077_lo_n
  );


  not

  (
    n1089_li,
    G40_n
  );


  not

  (
    n1092_li,
    n1089_lo_n
  );


  not

  (
    n1101_li,
    G41_n
  );


  not

  (
    n1104_li,
    n1101_lo_n
  );


  not

  (
    n1837_i2,
    n2151_o2_n_spl_
  );


  not

  (
    n1838_i2,
    n2152_o2_n_spl_
  );


  not

  (
    n1839_i2,
    n2153_o2_n_spl_
  );


  not

  (
    n1840_i2,
    n2154_o2_n_spl_
  );


  not

  (
    n1841_i2,
    n2155_o2_n_spl_
  );


  not

  (
    n1842_i2,
    n2156_o2_n_spl_
  );


  not

  (
    n1843_i2,
    n2157_o2_n_spl_
  );


  not

  (
    n1844_i2,
    n2158_o2_n_spl_
  );


  not

  (
    n1845_i2,
    n2159_o2_n_spl_
  );


  not

  (
    n1846_i2,
    n2160_o2_n_spl_
  );


  not

  (
    n1847_i2,
    n2161_o2_n_spl_
  );


  not

  (
    n1848_i2,
    n2162_o2_n_spl_
  );


  not

  (
    n1849_i2,
    n2163_o2_n_spl_
  );


  not

  (
    n1850_i2,
    n2164_o2_n_spl_
  );


  not

  (
    n1851_i2,
    n2165_o2_n_spl_
  );


  not

  (
    n1852_i2,
    n2166_o2_n_spl_
  );


  not

  (
    n1853_i2,
    n2167_o2_n_spl_
  );


  not

  (
    n1854_i2,
    n2168_o2_n_spl_
  );


  not

  (
    n1855_i2,
    n2169_o2_n_spl_
  );


  not

  (
    n1856_i2,
    n2170_o2_n_spl_
  );


  not

  (
    n1857_i2,
    n2171_o2_n_spl_
  );


  not

  (
    n1858_i2,
    n2172_o2_n_spl_
  );


  not

  (
    n1859_i2,
    n2173_o2_n_spl_
  );


  not

  (
    n1860_i2,
    n2174_o2_n_spl_
  );


  not

  (
    n1861_i2,
    n2175_o2_n_spl_
  );


  not

  (
    n1862_i2,
    n2176_o2_n_spl_
  );


  not

  (
    n1863_i2,
    n2177_o2_n_spl_
  );


  not

  (
    n1864_i2,
    n2178_o2_n_spl_
  );


  not

  (
    n1865_i2,
    n2179_o2_n_spl_
  );


  not

  (
    n1866_i2,
    n2180_o2_n_spl_
  );


  not

  (
    n1867_i2,
    n2181_o2_n_spl_
  );


  not

  (
    n1868_i2,
    n2182_o2_n_spl_
  );


  not

  (
    G834_i2,
    g433_p_spl_0
  );


  not

  (
    G847_i2,
    g437_p_spl_0
  );


  not

  (
    G860_i2,
    g441_p_spl_0
  );


  not

  (
    G873_i2,
    g445_p_spl_0
  );


  not

  (
    G925_i2,
    g449_p_spl_0
  );


  not

  (
    G886_i2,
    g453_p_spl_0
  );


  not

  (
    G912_i2,
    g457_p_spl_0
  );


  not

  (
    G899_i2,
    g461_p_spl_0
  );


  not

  (
    n2151_i2,
    n627_lo_buf_o2_n_spl_
  );


  not

  (
    n2152_i2,
    n639_lo_buf_o2_n_spl_
  );


  not

  (
    n2153_i2,
    n651_lo_buf_o2_n_spl_
  );


  not

  (
    n2154_i2,
    n663_lo_buf_o2_n_spl_
  );


  not

  (
    n2155_i2,
    n675_lo_buf_o2_n_spl_
  );


  not

  (
    n2156_i2,
    n687_lo_buf_o2_n_spl_
  );


  not

  (
    n2157_i2,
    n699_lo_buf_o2_n_spl_
  );


  not

  (
    n2158_i2,
    n711_lo_buf_o2_n_spl_
  );


  not

  (
    n2159_i2,
    n723_lo_buf_o2_n_spl_
  );


  not

  (
    n2160_i2,
    n735_lo_buf_o2_n_spl_
  );


  not

  (
    n2161_i2,
    n747_lo_buf_o2_n_spl_
  );


  not

  (
    n2162_i2,
    n759_lo_buf_o2_n_spl_
  );


  not

  (
    n2163_i2,
    n771_lo_buf_o2_n_spl_
  );


  not

  (
    n2164_i2,
    n783_lo_buf_o2_n_spl_
  );


  not

  (
    n2165_i2,
    n795_lo_buf_o2_n_spl_
  );


  not

  (
    n2166_i2,
    n807_lo_buf_o2_n_spl_
  );


  not

  (
    n2167_i2,
    n819_lo_buf_o2_n_spl_
  );


  not

  (
    n2168_i2,
    n831_lo_buf_o2_n_spl_
  );


  not

  (
    n2169_i2,
    n843_lo_buf_o2_n_spl_
  );


  not

  (
    n2170_i2,
    n855_lo_buf_o2_n_spl_
  );


  not

  (
    n2171_i2,
    n867_lo_buf_o2_n_spl_
  );


  not

  (
    n2172_i2,
    n879_lo_buf_o2_n_spl_
  );


  not

  (
    n2173_i2,
    n891_lo_buf_o2_n_spl_
  );


  not

  (
    n2174_i2,
    n903_lo_buf_o2_n_spl_
  );


  not

  (
    n2175_i2,
    n915_lo_buf_o2_n_spl_
  );


  not

  (
    n2176_i2,
    n927_lo_buf_o2_n_spl_
  );


  not

  (
    n2177_i2,
    n939_lo_buf_o2_n_spl_
  );


  not

  (
    n2178_i2,
    n951_lo_buf_o2_n_spl_
  );


  not

  (
    n2179_i2,
    n963_lo_buf_o2_n_spl_
  );


  not

  (
    n2180_i2,
    n975_lo_buf_o2_n_spl_
  );


  not

  (
    n2181_i2,
    n987_lo_buf_o2_n_spl_
  );


  not

  (
    n2182_i2,
    n999_lo_buf_o2_n_spl_
  );


  not

  (
    G974_i2,
    g433_p_spl_1
  );


  not

  (
    G976_i2,
    g433_p_spl_1
  );


  not

  (
    G970_i2,
    g437_p_spl_1
  );


  not

  (
    G972_i2,
    g437_p_spl_1
  );


  not

  (
    G973_i2,
    g441_p_spl_1
  );


  not

  (
    G977_i2,
    g441_p_spl_1
  );


  not

  (
    G971_i2,
    g445_p_spl_1
  );


  not

  (
    G975_i2,
    g445_p_spl_1
  );


  not

  (
    G954_i2,
    g449_p_spl_1
  );


  not

  (
    G956_i2,
    g449_p_spl_1
  );


  not

  (
    G950_i2,
    g453_p_spl_1
  );


  not

  (
    G952_i2,
    g453_p_spl_1
  );


  not

  (
    G953_i2,
    g457_p_spl_1
  );


  not

  (
    G957_i2,
    g457_p_spl_1
  );


  not

  (
    G951_i2,
    g461_p_spl_1
  );


  not

  (
    G955_i2,
    g461_p_spl_1
  );


  not

  (
    G986_i2,
    g475_p
  );


  not

  (
    G991_i2,
    g489_p
  );


  not

  (
    G770_i2,
    g498_p
  );


  not

  (
    G773_i2,
    g507_p
  );


  not

  (
    G776_i2,
    g516_p
  );


  not

  (
    G779_i2,
    g525_p
  );


  not

  (
    G782_i2,
    g534_p
  );


  not

  (
    G785_i2,
    g543_p
  );


  not

  (
    G788_i2,
    g552_p
  );


  not

  (
    G791_i2,
    g561_p
  );


  not

  (
    G642_i2,
    g573_p
  );


  not

  (
    G645_i2,
    g585_p
  );


  not

  (
    G648_i2,
    g597_p
  );


  not

  (
    G651_i2,
    g609_p
  );


  not

  (
    G654_i2,
    g621_p
  );


  not

  (
    G657_i2,
    g633_p
  );


  not

  (
    G660_i2,
    g645_p
  );


  not

  (
    G663_i2,
    g657_p
  );


  not

  (
    G602_i2,
    g669_p
  );


  not

  (
    G607_i2,
    g681_p
  );


  not

  (
    G612_i2,
    g693_p
  );


  not

  (
    G617_i2,
    g705_p
  );


  not

  (
    G622_i2,
    g717_p
  );


  not

  (
    G627_i2,
    g729_p
  );


  not

  (
    G632_i2,
    g741_p
  );


  not

  (
    G637_i2,
    g753_p
  );


  not

  (
    n627_lo_buf_i2,
    G1_n
  );


  not

  (
    n639_lo_buf_i2,
    G2_n
  );


  not

  (
    n651_lo_buf_i2,
    G3_n
  );


  not

  (
    n663_lo_buf_i2,
    G4_n
  );


  not

  (
    n675_lo_buf_i2,
    G5_n
  );


  not

  (
    n687_lo_buf_i2,
    G6_n
  );


  not

  (
    n699_lo_buf_i2,
    G7_n
  );


  not

  (
    n711_lo_buf_i2,
    G8_n
  );


  not

  (
    n723_lo_buf_i2,
    G9_n
  );


  not

  (
    n735_lo_buf_i2,
    G10_n
  );


  not

  (
    n747_lo_buf_i2,
    G11_n
  );


  not

  (
    n759_lo_buf_i2,
    G12_n
  );


  not

  (
    n771_lo_buf_i2,
    G13_n
  );


  not

  (
    n783_lo_buf_i2,
    G14_n
  );


  not

  (
    n795_lo_buf_i2,
    G15_n
  );


  not

  (
    n807_lo_buf_i2,
    G16_n
  );


  not

  (
    n819_lo_buf_i2,
    G17_n
  );


  not

  (
    n831_lo_buf_i2,
    G18_n
  );


  not

  (
    n843_lo_buf_i2,
    G19_n
  );


  not

  (
    n855_lo_buf_i2,
    G20_n
  );


  not

  (
    n867_lo_buf_i2,
    G21_n
  );


  not

  (
    n879_lo_buf_i2,
    G22_n
  );


  not

  (
    n891_lo_buf_i2,
    G23_n
  );


  not

  (
    n903_lo_buf_i2,
    G24_n
  );


  not

  (
    n915_lo_buf_i2,
    G25_n
  );


  not

  (
    n927_lo_buf_i2,
    G26_n
  );


  not

  (
    n939_lo_buf_i2,
    G27_n
  );


  not

  (
    n951_lo_buf_i2,
    G28_n
  );


  not

  (
    n963_lo_buf_i2,
    G29_n
  );


  not

  (
    n975_lo_buf_i2,
    G30_n
  );


  not

  (
    n987_lo_buf_i2,
    G31_n
  );


  not

  (
    n999_lo_buf_i2,
    G32_n
  );


  buf

  (
    G925_o2_p_spl_,
    G925_o2_p
  );


  buf

  (
    G925_o2_p_spl_0,
    G925_o2_p_spl_
  );


  buf

  (
    G925_o2_p_spl_00,
    G925_o2_p_spl_0
  );


  buf

  (
    G925_o2_p_spl_01,
    G925_o2_p_spl_0
  );


  buf

  (
    G925_o2_p_spl_1,
    G925_o2_p_spl_
  );


  buf

  (
    G925_o2_n_spl_,
    G925_o2_n
  );


  buf

  (
    G925_o2_n_spl_0,
    G925_o2_n_spl_
  );


  buf

  (
    G925_o2_n_spl_00,
    G925_o2_n_spl_0
  );


  buf

  (
    G925_o2_n_spl_01,
    G925_o2_n_spl_0
  );


  buf

  (
    G925_o2_n_spl_1,
    G925_o2_n_spl_
  );


  buf

  (
    G912_o2_p_spl_,
    G912_o2_p
  );


  buf

  (
    G912_o2_p_spl_0,
    G912_o2_p_spl_
  );


  buf

  (
    G912_o2_p_spl_00,
    G912_o2_p_spl_0
  );


  buf

  (
    G912_o2_p_spl_01,
    G912_o2_p_spl_0
  );


  buf

  (
    G912_o2_p_spl_1,
    G912_o2_p_spl_
  );


  buf

  (
    G912_o2_n_spl_,
    G912_o2_n
  );


  buf

  (
    G912_o2_n_spl_0,
    G912_o2_n_spl_
  );


  buf

  (
    G912_o2_n_spl_00,
    G912_o2_n_spl_0
  );


  buf

  (
    G912_o2_n_spl_01,
    G912_o2_n_spl_0
  );


  buf

  (
    G912_o2_n_spl_1,
    G912_o2_n_spl_
  );


  buf

  (
    G986_o2_p_spl_,
    G986_o2_p
  );


  buf

  (
    G986_o2_p_spl_0,
    G986_o2_p_spl_
  );


  buf

  (
    G986_o2_p_spl_1,
    G986_o2_p_spl_
  );


  buf

  (
    G986_o2_n_spl_,
    G986_o2_n
  );


  buf

  (
    G986_o2_n_spl_0,
    G986_o2_n_spl_
  );


  buf

  (
    G986_o2_n_spl_1,
    G986_o2_n_spl_
  );


  buf

  (
    g241_p_spl_,
    g241_p
  );


  buf

  (
    g241_p_spl_0,
    g241_p_spl_
  );


  buf

  (
    g241_p_spl_1,
    g241_p_spl_
  );


  buf

  (
    G834_o2_p_spl_,
    G834_o2_p
  );


  buf

  (
    G834_o2_p_spl_0,
    G834_o2_p_spl_
  );


  buf

  (
    G834_o2_p_spl_00,
    G834_o2_p_spl_0
  );


  buf

  (
    G834_o2_p_spl_01,
    G834_o2_p_spl_0
  );


  buf

  (
    G834_o2_p_spl_1,
    G834_o2_p_spl_
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    g241_n_spl_0,
    g241_n_spl_
  );


  buf

  (
    g241_n_spl_1,
    g241_n_spl_
  );


  buf

  (
    G834_o2_n_spl_,
    G834_o2_n
  );


  buf

  (
    G834_o2_n_spl_0,
    G834_o2_n_spl_
  );


  buf

  (
    G834_o2_n_spl_00,
    G834_o2_n_spl_0
  );


  buf

  (
    G834_o2_n_spl_01,
    G834_o2_n_spl_0
  );


  buf

  (
    G834_o2_n_spl_1,
    G834_o2_n_spl_
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    G847_o2_p_spl_,
    G847_o2_p
  );


  buf

  (
    G847_o2_p_spl_0,
    G847_o2_p_spl_
  );


  buf

  (
    G847_o2_p_spl_00,
    G847_o2_p_spl_0
  );


  buf

  (
    G847_o2_p_spl_01,
    G847_o2_p_spl_0
  );


  buf

  (
    G847_o2_p_spl_1,
    G847_o2_p_spl_
  );


  buf

  (
    G847_o2_n_spl_,
    G847_o2_n
  );


  buf

  (
    G847_o2_n_spl_0,
    G847_o2_n_spl_
  );


  buf

  (
    G847_o2_n_spl_00,
    G847_o2_n_spl_0
  );


  buf

  (
    G847_o2_n_spl_01,
    G847_o2_n_spl_0
  );


  buf

  (
    G847_o2_n_spl_1,
    G847_o2_n_spl_
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    G860_o2_p_spl_,
    G860_o2_p
  );


  buf

  (
    G860_o2_p_spl_0,
    G860_o2_p_spl_
  );


  buf

  (
    G860_o2_p_spl_00,
    G860_o2_p_spl_0
  );


  buf

  (
    G860_o2_p_spl_01,
    G860_o2_p_spl_0
  );


  buf

  (
    G860_o2_p_spl_1,
    G860_o2_p_spl_
  );


  buf

  (
    G860_o2_n_spl_,
    G860_o2_n
  );


  buf

  (
    G860_o2_n_spl_0,
    G860_o2_n_spl_
  );


  buf

  (
    G860_o2_n_spl_00,
    G860_o2_n_spl_0
  );


  buf

  (
    G860_o2_n_spl_01,
    G860_o2_n_spl_0
  );


  buf

  (
    G860_o2_n_spl_1,
    G860_o2_n_spl_
  );


  buf

  (
    g253_n_spl_,
    g253_n
  );


  buf

  (
    G873_o2_p_spl_,
    G873_o2_p
  );


  buf

  (
    G873_o2_p_spl_0,
    G873_o2_p_spl_
  );


  buf

  (
    G873_o2_p_spl_00,
    G873_o2_p_spl_0
  );


  buf

  (
    G873_o2_p_spl_01,
    G873_o2_p_spl_0
  );


  buf

  (
    G873_o2_p_spl_1,
    G873_o2_p_spl_
  );


  buf

  (
    G873_o2_n_spl_,
    G873_o2_n
  );


  buf

  (
    G873_o2_n_spl_0,
    G873_o2_n_spl_
  );


  buf

  (
    G873_o2_n_spl_00,
    G873_o2_n_spl_0
  );


  buf

  (
    G873_o2_n_spl_01,
    G873_o2_n_spl_0
  );


  buf

  (
    G873_o2_n_spl_1,
    G873_o2_n_spl_
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    G899_o2_p_spl_,
    G899_o2_p
  );


  buf

  (
    G899_o2_p_spl_0,
    G899_o2_p_spl_
  );


  buf

  (
    G899_o2_p_spl_00,
    G899_o2_p_spl_0
  );


  buf

  (
    G899_o2_p_spl_01,
    G899_o2_p_spl_0
  );


  buf

  (
    G899_o2_p_spl_1,
    G899_o2_p_spl_
  );


  buf

  (
    G899_o2_n_spl_,
    G899_o2_n
  );


  buf

  (
    G899_o2_n_spl_0,
    G899_o2_n_spl_
  );


  buf

  (
    G899_o2_n_spl_00,
    G899_o2_n_spl_0
  );


  buf

  (
    G899_o2_n_spl_01,
    G899_o2_n_spl_0
  );


  buf

  (
    G899_o2_n_spl_1,
    G899_o2_n_spl_
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g265_p_spl_0,
    g265_p_spl_
  );


  buf

  (
    g265_p_spl_1,
    g265_p_spl_
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g265_n_spl_0,
    g265_n_spl_
  );


  buf

  (
    g265_n_spl_1,
    g265_n_spl_
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    g282_n_spl_,
    g282_n
  );


  buf

  (
    G886_o2_p_spl_,
    G886_o2_p
  );


  buf

  (
    G886_o2_p_spl_0,
    G886_o2_p_spl_
  );


  buf

  (
    G886_o2_p_spl_00,
    G886_o2_p_spl_0
  );


  buf

  (
    G886_o2_p_spl_01,
    G886_o2_p_spl_0
  );


  buf

  (
    G886_o2_p_spl_1,
    G886_o2_p_spl_
  );


  buf

  (
    G886_o2_n_spl_,
    G886_o2_n
  );


  buf

  (
    G886_o2_n_spl_0,
    G886_o2_n_spl_
  );


  buf

  (
    G886_o2_n_spl_00,
    G886_o2_n_spl_0
  );


  buf

  (
    G886_o2_n_spl_01,
    G886_o2_n_spl_0
  );


  buf

  (
    G886_o2_n_spl_1,
    G886_o2_n_spl_
  );


  buf

  (
    g289_p_spl_,
    g289_p
  );


  buf

  (
    g289_p_spl_0,
    g289_p_spl_
  );


  buf

  (
    g289_p_spl_1,
    g289_p_spl_
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g289_n_spl_0,
    g289_n_spl_
  );


  buf

  (
    g289_n_spl_1,
    g289_n_spl_
  );


  buf

  (
    g291_n_spl_,
    g291_n
  );


  buf

  (
    g296_n_spl_,
    g296_n
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g306_n_spl_,
    g306_n
  );


  buf

  (
    g313_p_spl_,
    g313_p
  );


  buf

  (
    g313_p_spl_0,
    g313_p_spl_
  );


  buf

  (
    g313_p_spl_1,
    g313_p_spl_
  );


  buf

  (
    g313_n_spl_,
    g313_n
  );


  buf

  (
    g313_n_spl_0,
    g313_n_spl_
  );


  buf

  (
    g313_n_spl_1,
    g313_n_spl_
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g325_n_spl_,
    g325_n
  );


  buf

  (
    g330_n_spl_,
    g330_n
  );


  buf

  (
    G991_o2_p_spl_,
    G991_o2_p
  );


  buf

  (
    G991_o2_p_spl_0,
    G991_o2_p_spl_
  );


  buf

  (
    G991_o2_p_spl_1,
    G991_o2_p_spl_
  );


  buf

  (
    G991_o2_n_spl_,
    G991_o2_n
  );


  buf

  (
    G991_o2_n_spl_0,
    G991_o2_n_spl_
  );


  buf

  (
    G991_o2_n_spl_1,
    G991_o2_n_spl_
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g337_p_spl_0,
    g337_p_spl_
  );


  buf

  (
    g337_p_spl_1,
    g337_p_spl_
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g337_n_spl_0,
    g337_n_spl_
  );


  buf

  (
    g337_n_spl_1,
    g337_n_spl_
  );


  buf

  (
    g339_n_spl_,
    g339_n
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g354_n_spl_,
    g354_n
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g361_p_spl_0,
    g361_p_spl_
  );


  buf

  (
    g361_p_spl_1,
    g361_p_spl_
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g361_n_spl_0,
    g361_n_spl_
  );


  buf

  (
    g361_n_spl_1,
    g361_n_spl_
  );


  buf

  (
    g363_n_spl_,
    g363_n
  );


  buf

  (
    g368_n_spl_,
    g368_n
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_1,
    g385_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_1,
    g385_n_spl_
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g409_p_spl_1,
    g409_p_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g409_n_spl_1,
    g409_n_spl_
  );


  buf

  (
    g411_n_spl_,
    g411_n
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    G642_o2_p_spl_,
    G642_o2_p
  );


  buf

  (
    G770_o2_p_spl_,
    G770_o2_p
  );


  buf

  (
    G642_o2_n_spl_,
    G642_o2_n
  );


  buf

  (
    G770_o2_n_spl_,
    G770_o2_n
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    G645_o2_p_spl_,
    G645_o2_p
  );


  buf

  (
    G773_o2_p_spl_,
    G773_o2_p
  );


  buf

  (
    G645_o2_n_spl_,
    G645_o2_n
  );


  buf

  (
    G773_o2_n_spl_,
    G773_o2_n
  );


  buf

  (
    g434_n_spl_,
    g434_n
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    G648_o2_p_spl_,
    G648_o2_p
  );


  buf

  (
    G776_o2_p_spl_,
    G776_o2_p
  );


  buf

  (
    G648_o2_n_spl_,
    G648_o2_n
  );


  buf

  (
    G776_o2_n_spl_,
    G776_o2_n
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    G651_o2_p_spl_,
    G651_o2_p
  );


  buf

  (
    G779_o2_p_spl_,
    G779_o2_p
  );


  buf

  (
    G651_o2_n_spl_,
    G651_o2_n
  );


  buf

  (
    G779_o2_n_spl_,
    G779_o2_n
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    G654_o2_p_spl_,
    G654_o2_p
  );


  buf

  (
    G782_o2_p_spl_,
    G782_o2_p
  );


  buf

  (
    G654_o2_n_spl_,
    G654_o2_n
  );


  buf

  (
    G782_o2_n_spl_,
    G782_o2_n
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    G657_o2_p_spl_,
    G657_o2_p
  );


  buf

  (
    G785_o2_p_spl_,
    G785_o2_p
  );


  buf

  (
    G657_o2_n_spl_,
    G657_o2_n
  );


  buf

  (
    G785_o2_n_spl_,
    G785_o2_n
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    G660_o2_p_spl_,
    G660_o2_p
  );


  buf

  (
    G788_o2_p_spl_,
    G788_o2_p
  );


  buf

  (
    G660_o2_n_spl_,
    G660_o2_n
  );


  buf

  (
    G788_o2_n_spl_,
    G788_o2_n
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    G663_o2_p_spl_,
    G663_o2_p
  );


  buf

  (
    G791_o2_p_spl_,
    G791_o2_p
  );


  buf

  (
    G663_o2_n_spl_,
    G663_o2_n
  );


  buf

  (
    G791_o2_n_spl_,
    G791_o2_n
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g437_n_spl_,
    g437_n
  );


  buf

  (
    g433_n_spl_,
    g433_n
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g441_n_spl_0,
    g441_n_spl_
  );


  buf

  (
    g445_p_spl_,
    g445_p
  );


  buf

  (
    g445_p_spl_0,
    g445_p_spl_
  );


  buf

  (
    g445_p_spl_1,
    g445_p_spl_
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g441_p_spl_0,
    g441_p_spl_
  );


  buf

  (
    g441_p_spl_1,
    g441_p_spl_
  );


  buf

  (
    g445_n_spl_,
    g445_n
  );


  buf

  (
    g445_n_spl_0,
    g445_n_spl_
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g437_p_spl_0,
    g437_p_spl_
  );


  buf

  (
    g437_p_spl_1,
    g437_p_spl_
  );


  buf

  (
    g433_p_spl_,
    g433_p
  );


  buf

  (
    g433_p_spl_0,
    g433_p_spl_
  );


  buf

  (
    g433_p_spl_1,
    g433_p_spl_
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g457_n_spl_0,
    g457_n_spl_
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g461_p_spl_0,
    g461_p_spl_
  );


  buf

  (
    g461_p_spl_1,
    g461_p_spl_
  );


  buf

  (
    g457_p_spl_,
    g457_p
  );


  buf

  (
    g457_p_spl_0,
    g457_p_spl_
  );


  buf

  (
    g457_p_spl_1,
    g457_p_spl_
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g461_n_spl_0,
    g461_n_spl_
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g453_p_spl_0,
    g453_p_spl_
  );


  buf

  (
    g453_p_spl_1,
    g453_p_spl_
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g449_p_spl_0,
    g449_p_spl_
  );


  buf

  (
    g449_p_spl_1,
    g449_p_spl_
  );


  buf

  (
    n1104_lo_p_spl_,
    n1104_lo_p
  );


  buf

  (
    n1104_lo_p_spl_0,
    n1104_lo_p_spl_
  );


  buf

  (
    n1104_lo_p_spl_00,
    n1104_lo_p_spl_0
  );


  buf

  (
    n1104_lo_p_spl_01,
    n1104_lo_p_spl_0
  );


  buf

  (
    n1104_lo_p_spl_1,
    n1104_lo_p_spl_
  );


  buf

  (
    n1104_lo_p_spl_10,
    n1104_lo_p_spl_1
  );


  buf

  (
    n1104_lo_p_spl_11,
    n1104_lo_p_spl_1
  );


  buf

  (
    n1104_lo_n_spl_,
    n1104_lo_n
  );


  buf

  (
    n1104_lo_n_spl_0,
    n1104_lo_n_spl_
  );


  buf

  (
    n1104_lo_n_spl_00,
    n1104_lo_n_spl_0
  );


  buf

  (
    n1104_lo_n_spl_01,
    n1104_lo_n_spl_0
  );


  buf

  (
    n1104_lo_n_spl_1,
    n1104_lo_n_spl_
  );


  buf

  (
    n1104_lo_n_spl_10,
    n1104_lo_n_spl_1
  );


  buf

  (
    n1104_lo_n_spl_11,
    n1104_lo_n_spl_1
  );


  buf

  (
    G627_o2_p_spl_,
    G627_o2_p
  );


  buf

  (
    G627_o2_p_spl_0,
    G627_o2_p_spl_
  );


  buf

  (
    G627_o2_p_spl_1,
    G627_o2_p_spl_
  );


  buf

  (
    G622_o2_p_spl_,
    G622_o2_p
  );


  buf

  (
    G622_o2_p_spl_0,
    G622_o2_p_spl_
  );


  buf

  (
    G622_o2_p_spl_1,
    G622_o2_p_spl_
  );


  buf

  (
    G627_o2_n_spl_,
    G627_o2_n
  );


  buf

  (
    G627_o2_n_spl_0,
    G627_o2_n_spl_
  );


  buf

  (
    G627_o2_n_spl_1,
    G627_o2_n_spl_
  );


  buf

  (
    G622_o2_n_spl_,
    G622_o2_n
  );


  buf

  (
    G622_o2_n_spl_0,
    G622_o2_n_spl_
  );


  buf

  (
    G622_o2_n_spl_1,
    G622_o2_n_spl_
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g491_p_spl_,
    g491_p
  );


  buf

  (
    g495_p_spl_,
    g495_p
  );


  buf

  (
    G637_o2_p_spl_,
    G637_o2_p
  );


  buf

  (
    G637_o2_p_spl_0,
    G637_o2_p_spl_
  );


  buf

  (
    G637_o2_p_spl_1,
    G637_o2_p_spl_
  );


  buf

  (
    G632_o2_p_spl_,
    G632_o2_p
  );


  buf

  (
    G632_o2_p_spl_0,
    G632_o2_p_spl_
  );


  buf

  (
    G632_o2_p_spl_1,
    G632_o2_p_spl_
  );


  buf

  (
    G637_o2_n_spl_,
    G637_o2_n
  );


  buf

  (
    G637_o2_n_spl_0,
    G637_o2_n_spl_
  );


  buf

  (
    G637_o2_n_spl_1,
    G637_o2_n_spl_
  );


  buf

  (
    G632_o2_n_spl_,
    G632_o2_n
  );


  buf

  (
    G632_o2_n_spl_0,
    G632_o2_n_spl_
  );


  buf

  (
    G632_o2_n_spl_1,
    G632_o2_n_spl_
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    G607_o2_p_spl_,
    G607_o2_p
  );


  buf

  (
    G607_o2_p_spl_0,
    G607_o2_p_spl_
  );


  buf

  (
    G607_o2_p_spl_1,
    G607_o2_p_spl_
  );


  buf

  (
    G602_o2_p_spl_,
    G602_o2_p
  );


  buf

  (
    G602_o2_p_spl_0,
    G602_o2_p_spl_
  );


  buf

  (
    G602_o2_p_spl_1,
    G602_o2_p_spl_
  );


  buf

  (
    G607_o2_n_spl_,
    G607_o2_n
  );


  buf

  (
    G607_o2_n_spl_0,
    G607_o2_n_spl_
  );


  buf

  (
    G607_o2_n_spl_1,
    G607_o2_n_spl_
  );


  buf

  (
    G602_o2_n_spl_,
    G602_o2_n
  );


  buf

  (
    G602_o2_n_spl_0,
    G602_o2_n_spl_
  );


  buf

  (
    G602_o2_n_spl_1,
    G602_o2_n_spl_
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    G617_o2_p_spl_,
    G617_o2_p
  );


  buf

  (
    G617_o2_p_spl_0,
    G617_o2_p_spl_
  );


  buf

  (
    G617_o2_p_spl_1,
    G617_o2_p_spl_
  );


  buf

  (
    G612_o2_p_spl_,
    G612_o2_p
  );


  buf

  (
    G612_o2_p_spl_0,
    G612_o2_p_spl_
  );


  buf

  (
    G612_o2_p_spl_1,
    G612_o2_p_spl_
  );


  buf

  (
    G617_o2_n_spl_,
    G617_o2_n
  );


  buf

  (
    G617_o2_n_spl_0,
    G617_o2_n_spl_
  );


  buf

  (
    G617_o2_n_spl_1,
    G617_o2_n_spl_
  );


  buf

  (
    G612_o2_n_spl_,
    G612_o2_n
  );


  buf

  (
    G612_o2_n_spl_0,
    G612_o2_n_spl_
  );


  buf

  (
    G612_o2_n_spl_1,
    G612_o2_n_spl_
  );


  buf

  (
    g536_n_spl_,
    g536_n
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g558_p_spl_,
    g558_p
  );


  buf

  (
    n2155_o2_p_spl_,
    n2155_o2_p
  );


  buf

  (
    n2151_o2_p_spl_,
    n2151_o2_p
  );


  buf

  (
    n2155_o2_n_spl_,
    n2155_o2_n
  );


  buf

  (
    n2155_o2_n_spl_0,
    n2155_o2_n_spl_
  );


  buf

  (
    n2151_o2_n_spl_,
    n2151_o2_n
  );


  buf

  (
    n2151_o2_n_spl_0,
    n2151_o2_n_spl_
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    n2163_o2_p_spl_,
    n2163_o2_p
  );


  buf

  (
    n2159_o2_p_spl_,
    n2159_o2_p
  );


  buf

  (
    n2163_o2_n_spl_,
    n2163_o2_n
  );


  buf

  (
    n2163_o2_n_spl_0,
    n2163_o2_n_spl_
  );


  buf

  (
    n2159_o2_n_spl_,
    n2159_o2_n
  );


  buf

  (
    n2159_o2_n_spl_0,
    n2159_o2_n_spl_
  );


  buf

  (
    g566_n_spl_,
    g566_n
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g570_p_spl_,
    g570_p
  );


  buf

  (
    n2156_o2_p_spl_,
    n2156_o2_p
  );


  buf

  (
    n2152_o2_p_spl_,
    n2152_o2_p
  );


  buf

  (
    n2156_o2_n_spl_,
    n2156_o2_n
  );


  buf

  (
    n2156_o2_n_spl_0,
    n2156_o2_n_spl_
  );


  buf

  (
    n2152_o2_n_spl_,
    n2152_o2_n
  );


  buf

  (
    n2152_o2_n_spl_0,
    n2152_o2_n_spl_
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    n2164_o2_p_spl_,
    n2164_o2_p
  );


  buf

  (
    n2160_o2_p_spl_,
    n2160_o2_p
  );


  buf

  (
    n2164_o2_n_spl_,
    n2164_o2_n
  );


  buf

  (
    n2164_o2_n_spl_0,
    n2164_o2_n_spl_
  );


  buf

  (
    n2160_o2_n_spl_,
    n2160_o2_n
  );


  buf

  (
    n2160_o2_n_spl_0,
    n2160_o2_n_spl_
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g578_p_spl_,
    g578_p
  );


  buf

  (
    g582_p_spl_,
    g582_p
  );


  buf

  (
    n2157_o2_p_spl_,
    n2157_o2_p
  );


  buf

  (
    n2153_o2_p_spl_,
    n2153_o2_p
  );


  buf

  (
    n2157_o2_n_spl_,
    n2157_o2_n
  );


  buf

  (
    n2157_o2_n_spl_0,
    n2157_o2_n_spl_
  );


  buf

  (
    n2153_o2_n_spl_,
    n2153_o2_n
  );


  buf

  (
    n2153_o2_n_spl_0,
    n2153_o2_n_spl_
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    n2165_o2_p_spl_,
    n2165_o2_p
  );


  buf

  (
    n2161_o2_p_spl_,
    n2161_o2_p
  );


  buf

  (
    n2165_o2_n_spl_,
    n2165_o2_n
  );


  buf

  (
    n2165_o2_n_spl_0,
    n2165_o2_n_spl_
  );


  buf

  (
    n2161_o2_n_spl_,
    n2161_o2_n
  );


  buf

  (
    n2161_o2_n_spl_0,
    n2161_o2_n_spl_
  );


  buf

  (
    g590_n_spl_,
    g590_n
  );


  buf

  (
    g590_p_spl_,
    g590_p
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    n2158_o2_p_spl_,
    n2158_o2_p
  );


  buf

  (
    n2154_o2_p_spl_,
    n2154_o2_p
  );


  buf

  (
    n2158_o2_n_spl_,
    n2158_o2_n
  );


  buf

  (
    n2158_o2_n_spl_0,
    n2158_o2_n_spl_
  );


  buf

  (
    n2154_o2_n_spl_,
    n2154_o2_n
  );


  buf

  (
    n2154_o2_n_spl_0,
    n2154_o2_n_spl_
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    n2166_o2_p_spl_,
    n2166_o2_p
  );


  buf

  (
    n2162_o2_p_spl_,
    n2162_o2_p
  );


  buf

  (
    n2166_o2_n_spl_,
    n2166_o2_n
  );


  buf

  (
    n2166_o2_n_spl_0,
    n2166_o2_n_spl_
  );


  buf

  (
    n2162_o2_n_spl_,
    n2162_o2_n
  );


  buf

  (
    n2162_o2_n_spl_0,
    n2162_o2_n_spl_
  );


  buf

  (
    g602_n_spl_,
    g602_n
  );


  buf

  (
    g602_p_spl_,
    g602_p
  );


  buf

  (
    g606_p_spl_,
    g606_p
  );


  buf

  (
    n2171_o2_p_spl_,
    n2171_o2_p
  );


  buf

  (
    n2167_o2_p_spl_,
    n2167_o2_p
  );


  buf

  (
    n2171_o2_n_spl_,
    n2171_o2_n
  );


  buf

  (
    n2171_o2_n_spl_0,
    n2171_o2_n_spl_
  );


  buf

  (
    n2167_o2_n_spl_,
    n2167_o2_n
  );


  buf

  (
    n2167_o2_n_spl_0,
    n2167_o2_n_spl_
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g610_p_spl_,
    g610_p
  );


  buf

  (
    n2179_o2_p_spl_,
    n2179_o2_p
  );


  buf

  (
    n2175_o2_p_spl_,
    n2175_o2_p
  );


  buf

  (
    n2179_o2_n_spl_,
    n2179_o2_n
  );


  buf

  (
    n2179_o2_n_spl_0,
    n2179_o2_n_spl_
  );


  buf

  (
    n2175_o2_n_spl_,
    n2175_o2_n
  );


  buf

  (
    n2175_o2_n_spl_0,
    n2175_o2_n_spl_
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    g618_p_spl_,
    g618_p
  );


  buf

  (
    n2172_o2_p_spl_,
    n2172_o2_p
  );


  buf

  (
    n2168_o2_p_spl_,
    n2168_o2_p
  );


  buf

  (
    n2172_o2_n_spl_,
    n2172_o2_n
  );


  buf

  (
    n2172_o2_n_spl_0,
    n2172_o2_n_spl_
  );


  buf

  (
    n2168_o2_n_spl_,
    n2168_o2_n
  );


  buf

  (
    n2168_o2_n_spl_0,
    n2168_o2_n_spl_
  );


  buf

  (
    g622_n_spl_,
    g622_n
  );


  buf

  (
    g622_p_spl_,
    g622_p
  );


  buf

  (
    n2180_o2_p_spl_,
    n2180_o2_p
  );


  buf

  (
    n2176_o2_p_spl_,
    n2176_o2_p
  );


  buf

  (
    n2180_o2_n_spl_,
    n2180_o2_n
  );


  buf

  (
    n2180_o2_n_spl_0,
    n2180_o2_n_spl_
  );


  buf

  (
    n2176_o2_n_spl_,
    n2176_o2_n
  );


  buf

  (
    n2176_o2_n_spl_0,
    n2176_o2_n_spl_
  );


  buf

  (
    g626_n_spl_,
    g626_n
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    n2173_o2_p_spl_,
    n2173_o2_p
  );


  buf

  (
    n2169_o2_p_spl_,
    n2169_o2_p
  );


  buf

  (
    n2173_o2_n_spl_,
    n2173_o2_n
  );


  buf

  (
    n2173_o2_n_spl_0,
    n2173_o2_n_spl_
  );


  buf

  (
    n2169_o2_n_spl_,
    n2169_o2_n
  );


  buf

  (
    n2169_o2_n_spl_0,
    n2169_o2_n_spl_
  );


  buf

  (
    g634_n_spl_,
    g634_n
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    n2181_o2_p_spl_,
    n2181_o2_p
  );


  buf

  (
    n2177_o2_p_spl_,
    n2177_o2_p
  );


  buf

  (
    n2181_o2_n_spl_,
    n2181_o2_n
  );


  buf

  (
    n2181_o2_n_spl_0,
    n2181_o2_n_spl_
  );


  buf

  (
    n2177_o2_n_spl_,
    n2177_o2_n
  );


  buf

  (
    n2177_o2_n_spl_0,
    n2177_o2_n_spl_
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g642_p_spl_,
    g642_p
  );


  buf

  (
    n2174_o2_p_spl_,
    n2174_o2_p
  );


  buf

  (
    n2170_o2_p_spl_,
    n2170_o2_p
  );


  buf

  (
    n2174_o2_n_spl_,
    n2174_o2_n
  );


  buf

  (
    n2174_o2_n_spl_0,
    n2174_o2_n_spl_
  );


  buf

  (
    n2170_o2_n_spl_,
    n2170_o2_n
  );


  buf

  (
    n2170_o2_n_spl_0,
    n2170_o2_n_spl_
  );


  buf

  (
    g646_n_spl_,
    g646_n
  );


  buf

  (
    g646_p_spl_,
    g646_p
  );


  buf

  (
    n2182_o2_p_spl_,
    n2182_o2_p
  );


  buf

  (
    n2178_o2_p_spl_,
    n2178_o2_p
  );


  buf

  (
    n2182_o2_n_spl_,
    n2182_o2_n
  );


  buf

  (
    n2182_o2_n_spl_0,
    n2182_o2_n_spl_
  );


  buf

  (
    n2178_o2_n_spl_,
    n2178_o2_n
  );


  buf

  (
    n2178_o2_n_spl_0,
    n2178_o2_n_spl_
  );


  buf

  (
    g650_n_spl_,
    g650_n
  );


  buf

  (
    g650_p_spl_,
    g650_p
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    n639_lo_buf_o2_p_spl_,
    n639_lo_buf_o2_p
  );


  buf

  (
    n627_lo_buf_o2_p_spl_,
    n627_lo_buf_o2_p
  );


  buf

  (
    n639_lo_buf_o2_n_spl_,
    n639_lo_buf_o2_n
  );


  buf

  (
    n639_lo_buf_o2_n_spl_0,
    n639_lo_buf_o2_n_spl_
  );


  buf

  (
    n627_lo_buf_o2_n_spl_,
    n627_lo_buf_o2_n
  );


  buf

  (
    n627_lo_buf_o2_n_spl_0,
    n627_lo_buf_o2_n_spl_
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_p_spl_,
    g658_p
  );


  buf

  (
    n663_lo_buf_o2_p_spl_,
    n663_lo_buf_o2_p
  );


  buf

  (
    n651_lo_buf_o2_p_spl_,
    n651_lo_buf_o2_p
  );


  buf

  (
    n663_lo_buf_o2_n_spl_,
    n663_lo_buf_o2_n
  );


  buf

  (
    n663_lo_buf_o2_n_spl_0,
    n663_lo_buf_o2_n_spl_
  );


  buf

  (
    n651_lo_buf_o2_n_spl_,
    n651_lo_buf_o2_n
  );


  buf

  (
    n651_lo_buf_o2_n_spl_0,
    n651_lo_buf_o2_n_spl_
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    g662_p_spl_,
    g662_p
  );


  buf

  (
    g666_p_spl_,
    g666_p
  );


  buf

  (
    n687_lo_buf_o2_p_spl_,
    n687_lo_buf_o2_p
  );


  buf

  (
    n675_lo_buf_o2_p_spl_,
    n675_lo_buf_o2_p
  );


  buf

  (
    n687_lo_buf_o2_n_spl_,
    n687_lo_buf_o2_n
  );


  buf

  (
    n687_lo_buf_o2_n_spl_0,
    n687_lo_buf_o2_n_spl_
  );


  buf

  (
    n675_lo_buf_o2_n_spl_,
    n675_lo_buf_o2_n
  );


  buf

  (
    n675_lo_buf_o2_n_spl_0,
    n675_lo_buf_o2_n_spl_
  );


  buf

  (
    g670_n_spl_,
    g670_n
  );


  buf

  (
    g670_p_spl_,
    g670_p
  );


  buf

  (
    n711_lo_buf_o2_p_spl_,
    n711_lo_buf_o2_p
  );


  buf

  (
    n699_lo_buf_o2_p_spl_,
    n699_lo_buf_o2_p
  );


  buf

  (
    n711_lo_buf_o2_n_spl_,
    n711_lo_buf_o2_n
  );


  buf

  (
    n711_lo_buf_o2_n_spl_0,
    n711_lo_buf_o2_n_spl_
  );


  buf

  (
    n699_lo_buf_o2_n_spl_,
    n699_lo_buf_o2_n
  );


  buf

  (
    n699_lo_buf_o2_n_spl_0,
    n699_lo_buf_o2_n_spl_
  );


  buf

  (
    g674_n_spl_,
    g674_n
  );


  buf

  (
    g674_p_spl_,
    g674_p
  );


  buf

  (
    g678_p_spl_,
    g678_p
  );


  buf

  (
    n735_lo_buf_o2_p_spl_,
    n735_lo_buf_o2_p
  );


  buf

  (
    n723_lo_buf_o2_p_spl_,
    n723_lo_buf_o2_p
  );


  buf

  (
    n735_lo_buf_o2_n_spl_,
    n735_lo_buf_o2_n
  );


  buf

  (
    n735_lo_buf_o2_n_spl_0,
    n735_lo_buf_o2_n_spl_
  );


  buf

  (
    n723_lo_buf_o2_n_spl_,
    n723_lo_buf_o2_n
  );


  buf

  (
    n723_lo_buf_o2_n_spl_0,
    n723_lo_buf_o2_n_spl_
  );


  buf

  (
    g682_n_spl_,
    g682_n
  );


  buf

  (
    g682_p_spl_,
    g682_p
  );


  buf

  (
    n759_lo_buf_o2_p_spl_,
    n759_lo_buf_o2_p
  );


  buf

  (
    n747_lo_buf_o2_p_spl_,
    n747_lo_buf_o2_p
  );


  buf

  (
    n759_lo_buf_o2_n_spl_,
    n759_lo_buf_o2_n
  );


  buf

  (
    n759_lo_buf_o2_n_spl_0,
    n759_lo_buf_o2_n_spl_
  );


  buf

  (
    n747_lo_buf_o2_n_spl_,
    n747_lo_buf_o2_n
  );


  buf

  (
    n747_lo_buf_o2_n_spl_0,
    n747_lo_buf_o2_n_spl_
  );


  buf

  (
    g686_n_spl_,
    g686_n
  );


  buf

  (
    g686_p_spl_,
    g686_p
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    n783_lo_buf_o2_p_spl_,
    n783_lo_buf_o2_p
  );


  buf

  (
    n771_lo_buf_o2_p_spl_,
    n771_lo_buf_o2_p
  );


  buf

  (
    n783_lo_buf_o2_n_spl_,
    n783_lo_buf_o2_n
  );


  buf

  (
    n783_lo_buf_o2_n_spl_0,
    n783_lo_buf_o2_n_spl_
  );


  buf

  (
    n771_lo_buf_o2_n_spl_,
    n771_lo_buf_o2_n
  );


  buf

  (
    n771_lo_buf_o2_n_spl_0,
    n771_lo_buf_o2_n_spl_
  );


  buf

  (
    g694_n_spl_,
    g694_n
  );


  buf

  (
    g694_p_spl_,
    g694_p
  );


  buf

  (
    n807_lo_buf_o2_p_spl_,
    n807_lo_buf_o2_p
  );


  buf

  (
    n795_lo_buf_o2_p_spl_,
    n795_lo_buf_o2_p
  );


  buf

  (
    n807_lo_buf_o2_n_spl_,
    n807_lo_buf_o2_n
  );


  buf

  (
    n807_lo_buf_o2_n_spl_0,
    n807_lo_buf_o2_n_spl_
  );


  buf

  (
    n795_lo_buf_o2_n_spl_,
    n795_lo_buf_o2_n
  );


  buf

  (
    n795_lo_buf_o2_n_spl_0,
    n795_lo_buf_o2_n_spl_
  );


  buf

  (
    g698_n_spl_,
    g698_n
  );


  buf

  (
    g698_p_spl_,
    g698_p
  );


  buf

  (
    g702_p_spl_,
    g702_p
  );


  buf

  (
    n831_lo_buf_o2_p_spl_,
    n831_lo_buf_o2_p
  );


  buf

  (
    n819_lo_buf_o2_p_spl_,
    n819_lo_buf_o2_p
  );


  buf

  (
    n831_lo_buf_o2_n_spl_,
    n831_lo_buf_o2_n
  );


  buf

  (
    n831_lo_buf_o2_n_spl_0,
    n831_lo_buf_o2_n_spl_
  );


  buf

  (
    n819_lo_buf_o2_n_spl_,
    n819_lo_buf_o2_n
  );


  buf

  (
    n819_lo_buf_o2_n_spl_0,
    n819_lo_buf_o2_n_spl_
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    n855_lo_buf_o2_p_spl_,
    n855_lo_buf_o2_p
  );


  buf

  (
    n843_lo_buf_o2_p_spl_,
    n843_lo_buf_o2_p
  );


  buf

  (
    n855_lo_buf_o2_n_spl_,
    n855_lo_buf_o2_n
  );


  buf

  (
    n855_lo_buf_o2_n_spl_0,
    n855_lo_buf_o2_n_spl_
  );


  buf

  (
    n843_lo_buf_o2_n_spl_,
    n843_lo_buf_o2_n
  );


  buf

  (
    n843_lo_buf_o2_n_spl_0,
    n843_lo_buf_o2_n_spl_
  );


  buf

  (
    g710_n_spl_,
    g710_n
  );


  buf

  (
    g710_p_spl_,
    g710_p
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    n879_lo_buf_o2_p_spl_,
    n879_lo_buf_o2_p
  );


  buf

  (
    n867_lo_buf_o2_p_spl_,
    n867_lo_buf_o2_p
  );


  buf

  (
    n879_lo_buf_o2_n_spl_,
    n879_lo_buf_o2_n
  );


  buf

  (
    n879_lo_buf_o2_n_spl_0,
    n879_lo_buf_o2_n_spl_
  );


  buf

  (
    n867_lo_buf_o2_n_spl_,
    n867_lo_buf_o2_n
  );


  buf

  (
    n867_lo_buf_o2_n_spl_0,
    n867_lo_buf_o2_n_spl_
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


  buf

  (
    g718_p_spl_,
    g718_p
  );


  buf

  (
    n903_lo_buf_o2_p_spl_,
    n903_lo_buf_o2_p
  );


  buf

  (
    n891_lo_buf_o2_p_spl_,
    n891_lo_buf_o2_p
  );


  buf

  (
    n903_lo_buf_o2_n_spl_,
    n903_lo_buf_o2_n
  );


  buf

  (
    n903_lo_buf_o2_n_spl_0,
    n903_lo_buf_o2_n_spl_
  );


  buf

  (
    n891_lo_buf_o2_n_spl_,
    n891_lo_buf_o2_n
  );


  buf

  (
    n891_lo_buf_o2_n_spl_0,
    n891_lo_buf_o2_n_spl_
  );


  buf

  (
    g722_n_spl_,
    g722_n
  );


  buf

  (
    g722_p_spl_,
    g722_p
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    n927_lo_buf_o2_p_spl_,
    n927_lo_buf_o2_p
  );


  buf

  (
    n915_lo_buf_o2_p_spl_,
    n915_lo_buf_o2_p
  );


  buf

  (
    n927_lo_buf_o2_n_spl_,
    n927_lo_buf_o2_n
  );


  buf

  (
    n927_lo_buf_o2_n_spl_0,
    n927_lo_buf_o2_n_spl_
  );


  buf

  (
    n915_lo_buf_o2_n_spl_,
    n915_lo_buf_o2_n
  );


  buf

  (
    n915_lo_buf_o2_n_spl_0,
    n915_lo_buf_o2_n_spl_
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    n951_lo_buf_o2_p_spl_,
    n951_lo_buf_o2_p
  );


  buf

  (
    n939_lo_buf_o2_p_spl_,
    n939_lo_buf_o2_p
  );


  buf

  (
    n951_lo_buf_o2_n_spl_,
    n951_lo_buf_o2_n
  );


  buf

  (
    n951_lo_buf_o2_n_spl_0,
    n951_lo_buf_o2_n_spl_
  );


  buf

  (
    n939_lo_buf_o2_n_spl_,
    n939_lo_buf_o2_n
  );


  buf

  (
    n939_lo_buf_o2_n_spl_0,
    n939_lo_buf_o2_n_spl_
  );


  buf

  (
    g734_n_spl_,
    g734_n
  );


  buf

  (
    g734_p_spl_,
    g734_p
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    n975_lo_buf_o2_p_spl_,
    n975_lo_buf_o2_p
  );


  buf

  (
    n963_lo_buf_o2_p_spl_,
    n963_lo_buf_o2_p
  );


  buf

  (
    n975_lo_buf_o2_n_spl_,
    n975_lo_buf_o2_n
  );


  buf

  (
    n975_lo_buf_o2_n_spl_0,
    n975_lo_buf_o2_n_spl_
  );


  buf

  (
    n963_lo_buf_o2_n_spl_,
    n963_lo_buf_o2_n
  );


  buf

  (
    n963_lo_buf_o2_n_spl_0,
    n963_lo_buf_o2_n_spl_
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g742_p_spl_,
    g742_p
  );


  buf

  (
    n999_lo_buf_o2_p_spl_,
    n999_lo_buf_o2_p
  );


  buf

  (
    n987_lo_buf_o2_p_spl_,
    n987_lo_buf_o2_p
  );


  buf

  (
    n999_lo_buf_o2_n_spl_,
    n999_lo_buf_o2_n
  );


  buf

  (
    n999_lo_buf_o2_n_spl_0,
    n999_lo_buf_o2_n_spl_
  );


  buf

  (
    n987_lo_buf_o2_n_spl_,
    n987_lo_buf_o2_n
  );


  buf

  (
    n987_lo_buf_o2_n_spl_0,
    n987_lo_buf_o2_n_spl_
  );


  buf

  (
    g746_n_spl_,
    g746_n
  );


  buf

  (
    g746_p_spl_,
    g746_p
  );


  buf

  (
    g750_p_spl_,
    g750_p
  );


endmodule
