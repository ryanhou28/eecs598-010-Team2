// Benchmark "mymod" written by ABC on Sun Nov  5 22:49:20 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36,
    G426, G427, G428, G429, G430, G431, G432  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36;
  output G426, G427, G428, G429, G430, G431, G432;
  reg n229_lo, n253_lo, n256_lo, n259_lo, n262_lo, n277_lo, n301_lo,
    n304_lo, n307_lo, n310_lo, n325_lo, n349_lo, n352_lo, n355_lo, n358_lo,
    n373_lo, n397_lo, n400_lo, n403_lo, n406_lo, n421_lo, n445_lo, n448_lo,
    n451_lo, n454_lo, n469_lo, n493_lo, n496_lo, n499_lo, n502_lo, n517_lo,
    n520_lo, n541_lo, n544_lo, n547_lo, n550_lo, n565_lo, n589_lo, n592_lo,
    n595_lo, n598_lo, n613_lo, n625_lo, n628_lo, n631_lo, n634_lo, n852_o2,
    n853_o2, n955_o2, n956_o2, n531_o2, n549_o2, n537_o2, n540_o2, n546_o2,
    n534_o2, n552_o2, n543_o2, n961_o2, n223_inv, n555_o2, n1009_o2,
    n1010_o2, n1011_o2, n1012_o2, lo026_buf_o2, lo074_buf_o2, lo090_buf_o2,
    lo122_buf_o2, n510_o2, n498_o2, n516_o2, n507_o2, lo106_buf_o2,
    n519_o2, n1029_o2, n1041_o2, n1043_o2, n1045_o2, n558_o2, n563_o2,
    lo094_buf_o2, lo102_buf_o2, n522_o2, n298_inv, n486_o2, n304_inv,
    n564_o2, n528_o2, n492_o2, n530_o2, n548_o2, n536_o2, n539_o2,
    lo025_buf_o2, lo073_buf_o2, lo089_buf_o2, lo121_buf_o2, n509_o2,
    n513_o2, n501_o2, n504_o2, n495_o2, n497_o2, n515_o2, n506_o2,
    lo010_buf_o2, lo042_buf_o2, lo058_buf_o2, lo138_buf_o2, lo014_buf_o2,
    lo022_buf_o2, lo030_buf_o2, lo038_buf_o2, lo046_buf_o2, lo054_buf_o2,
    lo126_buf_o2, lo134_buf_o2, lo093_buf_o2, lo101_buf_o2, lo002_buf_o2,
    lo006_buf_o2, lo062_buf_o2, lo070_buf_o2, lo078_buf_o2, lo086_buf_o2,
    lo110_buf_o2, lo118_buf_o2, n476_o2, n482_o2, n478_o2, n479_o2;
  wire new_n308_, new_n310_, new_n312_, new_n314_, new_n315_, new_n316_,
    new_n318_, new_n320_, new_n322_, new_n323_, new_n324_, new_n326_,
    new_n328_, new_n330_, new_n331_, new_n332_, new_n334_, new_n336_,
    new_n338_, new_n340_, new_n342_, new_n344_, new_n346_, new_n348_,
    new_n350_, new_n352_, new_n354_, new_n356_, new_n358_, new_n360_,
    new_n362_, new_n364_, new_n366_, new_n368_, new_n370_, new_n371_,
    new_n372_, new_n374_, new_n376_, new_n378_, new_n380_, new_n382_,
    new_n384_, new_n386_, new_n389_, new_n390_, new_n392_, new_n394_,
    new_n396_, new_n398_, new_n400_, new_n402_, new_n404_, new_n406_,
    new_n408_, new_n409_, new_n410_, new_n412_, new_n414_, new_n416_,
    new_n418_, new_n419_, new_n420_, new_n422_, new_n424_, new_n426_,
    new_n428_, new_n429_, new_n430_, new_n432_, new_n434_, new_n436_,
    new_n438_, new_n440_, new_n442_, new_n444_, new_n446_, new_n448_,
    new_n450_, new_n451_, new_n452_, new_n454_, new_n456_, new_n458_,
    new_n460_, new_n462_, new_n464_, new_n466_, new_n468_, new_n470_,
    new_n472_, new_n474_, new_n476_, new_n478_, new_n480_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n487_, new_n489_, new_n490_,
    new_n491_, new_n493_, new_n495_, new_n496_, new_n498_, new_n500_,
    new_n501_, new_n503_, new_n505_, new_n507_, new_n509_, new_n510_,
    new_n512_, new_n514_, new_n516_, new_n519_, new_n521_, new_n523_,
    new_n525_, new_n526_, new_n529_, new_n531_, new_n533_, new_n535_,
    new_n537_, new_n538_, new_n540_, new_n542_, new_n545_, new_n546_,
    new_n548_, new_n550_, new_n552_, new_n554_, new_n555_, new_n556_,
    new_n558_, new_n560_, new_n562_, new_n564_, new_n566_, new_n568_,
    new_n570_, new_n572_, new_n574_, new_n576_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n604_, new_n607_, new_n608_, new_n611_, new_n612_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n638_, new_n640_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, n856_li008_li008, n880_li016_li016,
    n883_li017_li017, n886_li018_li018, n889_li019_li019, n904_li024_li024,
    n928_li032_li032, n931_li033_li033, n934_li034_li034, n937_li035_li035,
    n952_li040_li040, n976_li048_li048, n979_li049_li049, n982_li050_li050,
    n985_li051_li051, n1000_li056_li056, n1024_li064_li064,
    n1027_li065_li065, n1030_li066_li066, n1033_li067_li067,
    n1048_li072_li072, n1072_li080_li080, n1075_li081_li081,
    n1078_li082_li082, n1081_li083_li083, n1096_li088_li088,
    n1120_li096_li096, n1123_li097_li097, n1126_li098_li098,
    n1129_li099_li099, n1144_li104_li104, n1147_li105_li105,
    n1168_li112_li112, n1171_li113_li113, n1174_li114_li114,
    n1177_li115_li115, n1192_li120_li120, n1216_li128_li128,
    n1219_li129_li129, n1222_li130_li130, n1225_li131_li131,
    n1240_li136_li136, n1252_li140_li140, n1255_li141_li141,
    n1258_li142_li142, n1261_li143_li143, n852_i2, n853_i2, n955_i2,
    n956_i2, n531_i2, n549_i2, n537_i2, n540_i2, n546_i2, n534_i2, n552_i2,
    n543_i2, n961_i2, n962_i2, n555_i2, n1009_i2, n1010_i2, n1011_i2,
    n1012_i2, lo026_buf_i2, lo074_buf_i2, lo090_buf_i2, lo122_buf_i2,
    n510_i2, n498_i2, n516_i2, n507_i2, lo106_buf_i2, n519_i2, n1029_i2,
    n1041_i2, n1043_i2, n1045_i2, n558_i2, n563_i2, lo094_buf_i2,
    lo102_buf_i2, n522_i2, n527_i2, n486_i2, n491_i2, n564_i2, n528_i2,
    n492_i2, n530_i2, n548_i2, n536_i2, n539_i2, lo025_buf_i2,
    lo073_buf_i2, lo089_buf_i2, lo121_buf_i2, n509_i2, n513_i2, n501_i2,
    n504_i2, n495_i2, n497_i2, n515_i2, n506_i2, lo010_buf_i2,
    lo042_buf_i2, lo058_buf_i2, lo138_buf_i2, lo014_buf_i2, lo022_buf_i2,
    lo030_buf_i2, lo038_buf_i2, lo046_buf_i2, lo054_buf_i2, lo126_buf_i2,
    lo134_buf_i2, lo093_buf_i2, lo101_buf_i2, lo002_buf_i2, lo006_buf_i2,
    lo062_buf_i2, lo070_buf_i2, lo078_buf_i2, lo086_buf_i2, lo110_buf_i2,
    lo118_buf_i2, n476_i2, n482_i2, n478_i2, n479_i2;
  assign new_n308_ = G1;
  assign new_n310_ = G2;
  assign new_n312_ = G3;
  assign new_n314_ = G4;
  assign new_n315_ = ~G4;
  assign new_n316_ = G5;
  assign new_n318_ = G6;
  assign new_n320_ = G7;
  assign new_n322_ = G8;
  assign new_n323_ = ~G8;
  assign new_n324_ = G9;
  assign new_n326_ = G10;
  assign new_n328_ = G11;
  assign new_n330_ = G12;
  assign new_n331_ = ~G12;
  assign new_n332_ = G13;
  assign new_n334_ = G14;
  assign new_n336_ = G15;
  assign new_n338_ = G16;
  assign new_n340_ = G17;
  assign new_n342_ = G18;
  assign new_n344_ = G19;
  assign new_n346_ = G20;
  assign new_n348_ = G21;
  assign new_n350_ = G22;
  assign new_n352_ = G23;
  assign new_n354_ = G24;
  assign new_n356_ = G25;
  assign new_n358_ = G26;
  assign new_n360_ = G27;
  assign new_n362_ = G28;
  assign new_n364_ = G29;
  assign new_n366_ = G30;
  assign new_n368_ = G31;
  assign new_n370_ = G32;
  assign new_n371_ = ~G32;
  assign new_n372_ = G33;
  assign new_n374_ = G34;
  assign new_n376_ = G35;
  assign new_n378_ = G36;
  assign new_n380_ = n229_lo;
  assign new_n382_ = n253_lo;
  assign new_n384_ = n256_lo;
  assign new_n386_ = n259_lo;
  assign new_n389_ = ~n262_lo;
  assign new_n390_ = n277_lo;
  assign new_n392_ = n301_lo;
  assign new_n394_ = n304_lo;
  assign new_n396_ = n307_lo;
  assign new_n398_ = n310_lo;
  assign new_n400_ = n325_lo;
  assign new_n402_ = n349_lo;
  assign new_n404_ = n352_lo;
  assign new_n406_ = n355_lo;
  assign new_n408_ = n358_lo;
  assign new_n409_ = ~n358_lo;
  assign new_n410_ = n373_lo;
  assign new_n412_ = n397_lo;
  assign new_n414_ = n400_lo;
  assign new_n416_ = n403_lo;
  assign new_n418_ = n406_lo;
  assign new_n419_ = ~n406_lo;
  assign new_n420_ = n421_lo;
  assign new_n422_ = n445_lo;
  assign new_n424_ = n448_lo;
  assign new_n426_ = n451_lo;
  assign new_n428_ = n454_lo;
  assign new_n429_ = ~n454_lo;
  assign new_n430_ = n469_lo;
  assign new_n432_ = n493_lo;
  assign new_n434_ = n496_lo;
  assign new_n436_ = n499_lo;
  assign new_n438_ = n502_lo;
  assign new_n440_ = n517_lo;
  assign new_n442_ = n520_lo;
  assign new_n444_ = n541_lo;
  assign new_n446_ = n544_lo;
  assign new_n448_ = n547_lo;
  assign new_n450_ = n550_lo;
  assign new_n451_ = ~n550_lo;
  assign new_n452_ = n565_lo;
  assign new_n454_ = n589_lo;
  assign new_n456_ = n592_lo;
  assign new_n458_ = n595_lo;
  assign new_n460_ = n598_lo;
  assign new_n462_ = n613_lo;
  assign new_n464_ = n625_lo;
  assign new_n466_ = n628_lo;
  assign new_n468_ = n631_lo;
  assign new_n470_ = n634_lo;
  assign new_n472_ = n852_o2;
  assign new_n474_ = n853_o2;
  assign new_n476_ = n955_o2;
  assign new_n478_ = n956_o2;
  assign new_n480_ = n531_o2;
  assign new_n482_ = n549_o2;
  assign new_n483_ = ~n549_o2;
  assign new_n484_ = n537_o2;
  assign new_n485_ = ~n537_o2;
  assign new_n487_ = ~n540_o2;
  assign new_n489_ = ~n546_o2;
  assign new_n490_ = n534_o2;
  assign new_n491_ = ~n534_o2;
  assign new_n493_ = ~n552_o2;
  assign new_n495_ = ~n543_o2;
  assign new_n496_ = n961_o2;
  assign new_n498_ = n223_inv;
  assign new_n500_ = n555_o2;
  assign new_n501_ = ~n555_o2;
  assign new_n503_ = ~n1009_o2;
  assign new_n505_ = ~n1010_o2;
  assign new_n507_ = ~n1011_o2;
  assign new_n509_ = ~n1012_o2;
  assign new_n510_ = lo026_buf_o2;
  assign new_n512_ = lo074_buf_o2;
  assign new_n514_ = lo090_buf_o2;
  assign new_n516_ = lo122_buf_o2;
  assign new_n519_ = ~n510_o2;
  assign new_n521_ = ~n498_o2;
  assign new_n523_ = ~n516_o2;
  assign new_n525_ = ~n507_o2;
  assign new_n526_ = lo106_buf_o2;
  assign new_n529_ = ~n519_o2;
  assign new_n531_ = ~n1029_o2;
  assign new_n533_ = ~n1041_o2;
  assign new_n535_ = ~n1043_o2;
  assign new_n537_ = ~n1045_o2;
  assign new_n538_ = n558_o2;
  assign new_n540_ = n563_o2;
  assign new_n542_ = lo094_buf_o2;
  assign new_n545_ = ~lo102_buf_o2;
  assign new_n546_ = n522_o2;
  assign new_n548_ = n298_inv;
  assign new_n550_ = n486_o2;
  assign new_n552_ = n304_inv;
  assign new_n554_ = n564_o2;
  assign new_n555_ = ~n564_o2;
  assign new_n556_ = n528_o2;
  assign new_n558_ = n492_o2;
  assign new_n560_ = n530_o2;
  assign new_n562_ = n548_o2;
  assign new_n564_ = n536_o2;
  assign new_n566_ = n539_o2;
  assign new_n568_ = lo025_buf_o2;
  assign new_n570_ = lo073_buf_o2;
  assign new_n572_ = lo089_buf_o2;
  assign new_n574_ = lo121_buf_o2;
  assign new_n576_ = n509_o2;
  assign new_n578_ = n513_o2;
  assign new_n579_ = ~n513_o2;
  assign new_n580_ = n501_o2;
  assign new_n581_ = ~n501_o2;
  assign new_n582_ = n504_o2;
  assign new_n583_ = ~n504_o2;
  assign new_n584_ = n495_o2;
  assign new_n585_ = ~n495_o2;
  assign new_n586_ = n497_o2;
  assign new_n588_ = n515_o2;
  assign new_n590_ = n506_o2;
  assign new_n592_ = lo010_buf_o2;
  assign new_n593_ = ~lo010_buf_o2;
  assign new_n594_ = lo042_buf_o2;
  assign new_n595_ = ~lo042_buf_o2;
  assign new_n596_ = lo058_buf_o2;
  assign new_n597_ = ~lo058_buf_o2;
  assign new_n598_ = lo138_buf_o2;
  assign new_n599_ = ~lo138_buf_o2;
  assign new_n600_ = lo014_buf_o2;
  assign new_n602_ = lo022_buf_o2;
  assign new_n604_ = lo030_buf_o2;
  assign new_n607_ = ~lo038_buf_o2;
  assign new_n608_ = lo046_buf_o2;
  assign new_n611_ = ~lo054_buf_o2;
  assign new_n612_ = lo126_buf_o2;
  assign new_n615_ = ~lo134_buf_o2;
  assign new_n616_ = lo093_buf_o2;
  assign new_n617_ = ~lo093_buf_o2;
  assign new_n618_ = lo101_buf_o2;
  assign new_n620_ = lo002_buf_o2;
  assign new_n621_ = ~lo002_buf_o2;
  assign new_n622_ = lo006_buf_o2;
  assign new_n623_ = ~lo006_buf_o2;
  assign new_n624_ = lo062_buf_o2;
  assign new_n625_ = ~lo062_buf_o2;
  assign new_n626_ = lo070_buf_o2;
  assign new_n628_ = lo078_buf_o2;
  assign new_n629_ = ~lo078_buf_o2;
  assign new_n630_ = lo086_buf_o2;
  assign new_n632_ = lo110_buf_o2;
  assign new_n633_ = ~lo110_buf_o2;
  assign new_n634_ = lo118_buf_o2;
  assign new_n636_ = n476_o2;
  assign new_n638_ = n482_o2;
  assign new_n640_ = n478_o2;
  assign new_n642_ = n479_o2;
  assign new_n644_ = new_n472_ | new_n474_;
  assign new_n645_ = new_n476_ | new_n478_;
  assign new_n646_ = new_n538_ | new_n540_;
  assign new_n647_ = new_n389_ | new_n921_;
  assign new_n648_ = new_n480_ & new_n647_;
  assign new_n649_ = new_n460_ & new_n925_;
  assign new_n650_ = new_n495_ | new_n649_;
  assign new_n651_ = new_n450_ & new_n925_;
  assign new_n652_ = new_n451_ | new_n921_;
  assign new_n653_ = new_n500_ & new_n652_;
  assign new_n654_ = new_n501_ | new_n651_;
  assign new_n655_ = new_n930_ & new_n931_;
  assign new_n656_ = new_n438_ & new_n926_;
  assign new_n657_ = new_n493_ | new_n656_;
  assign new_n658_ = new_n470_ & new_n926_;
  assign new_n659_ = new_n487_ | new_n658_;
  assign new_n660_ = new_n932_ & new_n659_;
  assign new_n661_ = new_n655_ & new_n660_;
  assign new_n662_ = new_n408_ & new_n928_;
  assign new_n663_ = new_n409_ | new_n920_;
  assign new_n664_ = new_n482_ & new_n663_;
  assign new_n665_ = new_n483_ | new_n662_;
  assign new_n666_ = new_n428_ & new_n928_;
  assign new_n667_ = new_n429_ | new_n922_;
  assign new_n668_ = new_n490_ & new_n667_;
  assign new_n669_ = new_n491_ | new_n666_;
  assign new_n670_ = new_n933_ & new_n669_;
  assign new_n671_ = new_n934_ | new_n935_;
  assign new_n672_ = new_n398_ & new_n929_;
  assign new_n673_ = new_n489_ | new_n672_;
  assign new_n674_ = new_n418_ & new_n929_;
  assign new_n675_ = new_n419_ | new_n922_;
  assign new_n676_ = new_n484_ & new_n675_;
  assign new_n677_ = new_n485_ | new_n674_;
  assign new_n678_ = new_n936_ & new_n937_;
  assign new_n679_ = new_n670_ & new_n678_;
  assign new_n680_ = new_n661_ & new_n938_;
  assign new_n681_ = new_n648_ | new_n680_;
  assign new_n682_ = new_n932_ | new_n939_;
  assign new_n683_ = new_n671_ | new_n682_;
  assign new_n684_ = new_n936_ & new_n683_;
  assign new_n685_ = new_n935_ | new_n939_;
  assign new_n686_ = new_n931_ | new_n685_;
  assign new_n687_ = new_n933_ & new_n686_;
  assign new_n688_ = new_n940_ & new_n687_;
  assign new_n689_ = new_n930_ | new_n653_;
  assign new_n690_ = new_n937_ & new_n689_;
  assign new_n691_ = new_n934_ | new_n690_;
  assign new_n692_ = new_n940_ & new_n691_;
  assign new_n693_ = new_n509_ | new_n560_;
  assign new_n694_ = new_n503_ | new_n562_;
  assign new_n695_ = new_n505_ | new_n564_;
  assign new_n696_ = new_n507_ | new_n566_;
  assign new_n697_ = new_n510_ & new_n943_;
  assign new_n698_ = new_n519_ | new_n697_;
  assign new_n699_ = new_n512_ & new_n943_;
  assign new_n700_ = new_n521_ | new_n699_;
  assign new_n701_ = new_n514_ & new_n942_;
  assign new_n702_ = new_n523_ | new_n701_;
  assign new_n703_ = new_n516_ & new_n944_;
  assign new_n704_ = new_n525_ | new_n703_;
  assign new_n705_ = new_n526_ & new_n944_;
  assign new_n706_ = new_n529_ | new_n705_;
  assign new_n707_ = new_n531_ | new_n576_;
  assign new_n708_ = new_n533_ | new_n586_;
  assign new_n709_ = new_n535_ | new_n588_;
  assign new_n710_ = new_n537_ | new_n590_;
  assign new_n711_ = new_n542_ & new_n558_;
  assign new_n712_ = new_n545_ | new_n711_;
  assign new_n713_ = new_n945_ | new_n946_;
  assign new_n714_ = new_n947_ | new_n948_;
  assign new_n715_ = new_n949_ | new_n950_;
  assign new_n716_ = new_n714_ & new_n715_;
  assign new_n717_ = new_n713_ & new_n716_;
  assign new_n718_ = new_n951_ | new_n952_;
  assign new_n719_ = new_n953_ | new_n954_;
  assign new_n720_ = new_n718_ & new_n719_;
  assign new_n721_ = new_n955_ | new_n956_;
  assign new_n722_ = new_n957_ | new_n958_;
  assign new_n723_ = new_n721_ & new_n722_;
  assign new_n724_ = new_n959_ | new_n960_;
  assign new_n725_ = new_n961_ | new_n962_;
  assign new_n726_ = new_n724_ & new_n725_;
  assign new_n727_ = new_n723_ & new_n726_;
  assign new_n728_ = new_n720_ & new_n727_;
  assign new_n729_ = new_n963_ | new_n964_;
  assign new_n730_ = new_n965_ | new_n966_;
  assign new_n731_ = new_n967_ | new_n968_;
  assign new_n732_ = new_n730_ & new_n731_;
  assign new_n733_ = new_n729_ & new_n732_;
  assign new_n734_ = new_n969_ | new_n970_;
  assign new_n735_ = new_n971_ | new_n972_;
  assign new_n736_ = new_n734_ & new_n735_;
  assign new_n737_ = new_n585_ | new_n592_;
  assign new_n738_ = new_n583_ | new_n598_;
  assign new_n739_ = new_n737_ & new_n738_;
  assign new_n740_ = new_n581_ | new_n596_;
  assign new_n741_ = new_n579_ | new_n594_;
  assign new_n742_ = new_n740_ & new_n741_;
  assign new_n743_ = new_n739_ & new_n742_;
  assign new_n744_ = new_n736_ & new_n743_;
  assign new_n745_ = new_n617_ & new_n973_;
  assign new_n746_ = new_n633_ & new_n974_;
  assign new_n747_ = new_n621_ & new_n622_;
  assign new_n748_ = new_n746_ | new_n747_;
  assign new_n749_ = new_n745_ | new_n748_;
  assign new_n750_ = new_n625_ & new_n975_;
  assign new_n751_ = new_n629_ & new_n976_;
  assign new_n752_ = new_n750_ | new_n751_;
  assign new_n753_ = new_n636_ | new_n642_;
  assign new_n754_ = new_n638_ | new_n640_;
  assign new_n755_ = new_n753_ | new_n754_;
  assign new_n756_ = new_n752_ | new_n755_;
  assign new_n757_ = new_n977_ & new_n978_;
  assign new_n758_ = new_n979_ & new_n980_;
  assign new_n759_ = new_n981_ | new_n982_;
  assign new_n760_ = new_n593_ | new_n985_;
  assign new_n761_ = new_n595_ | new_n985_;
  assign new_n762_ = new_n597_ | new_n984_;
  assign new_n763_ = new_n599_ | new_n986_;
  assign new_n764_ = new_n600_ & new_n990_;
  assign new_n765_ = new_n604_ & new_n990_;
  assign new_n766_ = new_n607_ | new_n765_;
  assign new_n767_ = new_n608_ & new_n989_;
  assign new_n768_ = new_n611_ | new_n767_;
  assign new_n769_ = new_n612_ & new_n991_;
  assign new_n770_ = new_n615_ | new_n769_;
  assign new_n771_ = new_n620_ & new_n991_;
  assign new_n772_ = new_n623_ | new_n771_;
  assign new_n773_ = new_n624_ & new_n993_;
  assign new_n774_ = new_n628_ & new_n993_;
  assign new_n775_ = new_n632_ & new_n994_;
  assign new_n776_ = new_n315_ & new_n995_;
  assign new_n777_ = new_n323_ & new_n996_;
  assign new_n778_ = new_n331_ & new_n997_;
  assign new_n779_ = new_n371_ & new_n998_;
  assign G426 = new_n644_;
  assign G427 = new_n645_;
  assign G428 = new_n646_;
  assign G429 = ~new_n681_;
  assign G430 = ~new_n938_;
  assign G431 = ~new_n688_;
  assign G432 = ~new_n692_;
  assign n856_li008_li008 = new_n312_;
  assign n880_li016_li016 = new_n316_;
  assign n883_li017_li017 = new_n382_;
  assign n886_li018_li018 = new_n384_;
  assign n889_li019_li019 = new_n955_;
  assign n904_li024_li024 = new_n320_;
  assign n928_li032_li032 = new_n324_;
  assign n931_li033_li033 = new_n392_;
  assign n934_li034_li034 = new_n394_;
  assign n937_li035_li035 = new_n949_;
  assign n952_li040_li040 = new_n328_;
  assign n976_li048_li048 = new_n332_;
  assign n979_li049_li049 = new_n402_;
  assign n982_li050_li050 = new_n404_;
  assign n985_li051_li051 = new_n961_;
  assign n1000_li056_li056 = new_n336_;
  assign n1024_li064_li064 = new_n340_;
  assign n1027_li065_li065 = new_n412_;
  assign n1030_li066_li066 = new_n414_;
  assign n1033_li067_li067 = new_n959_;
  assign n1048_li072_li072 = new_n344_;
  assign n1072_li080_li080 = new_n348_;
  assign n1075_li081_li081 = new_n422_;
  assign n1078_li082_li082 = new_n424_;
  assign n1081_li083_li083 = new_n951_;
  assign n1096_li088_li088 = new_n352_;
  assign n1120_li096_li096 = new_n356_;
  assign n1123_li097_li097 = new_n432_;
  assign n1126_li098_li098 = new_n434_;
  assign n1129_li099_li099 = new_n953_;
  assign n1144_li104_li104 = new_n360_;
  assign n1147_li105_li105 = new_n440_;
  assign n1168_li112_li112 = new_n364_;
  assign n1171_li113_li113 = new_n444_;
  assign n1174_li114_li114 = new_n446_;
  assign n1177_li115_li115 = new_n945_;
  assign n1192_li120_li120 = new_n368_;
  assign n1216_li128_li128 = new_n372_;
  assign n1219_li129_li129 = new_n454_;
  assign n1222_li130_li130 = new_n456_;
  assign n1225_li131_li131 = new_n947_;
  assign n1240_li136_li136 = new_n376_;
  assign n1252_li140_li140 = new_n378_;
  assign n1255_li141_li141 = new_n464_;
  assign n1258_li142_li142 = new_n466_;
  assign n1261_li143_li143 = new_n957_;
  assign n852_i2 = new_n496_;
  assign n853_i2 = new_n498_;
  assign n955_i2 = new_n546_;
  assign n956_i2 = new_n548_;
  assign n531_i2 = ~new_n956_;
  assign n549_i2 = ~new_n962_;
  assign n537_i2 = ~new_n960_;
  assign n540_i2 = ~new_n958_;
  assign n546_i2 = ~new_n950_;
  assign n534_i2 = ~new_n952_;
  assign n552_i2 = ~new_n954_;
  assign n543_i2 = ~new_n948_;
  assign n961_i2 = new_n550_;
  assign n962_i2 = new_n552_;
  assign n555_i2 = ~new_n946_;
  assign n1009_i2 = new_n578_;
  assign n1010_i2 = new_n580_;
  assign n1011_i2 = new_n582_;
  assign n1012_i2 = new_n584_;
  assign lo026_buf_i2 = new_n967_;
  assign lo074_buf_i2 = new_n969_;
  assign lo090_buf_i2 = new_n971_;
  assign lo122_buf_i2 = new_n965_;
  assign n510_i2 = ~new_n968_;
  assign n498_i2 = ~new_n970_;
  assign n516_i2 = ~new_n972_;
  assign n507_i2 = ~new_n966_;
  assign lo106_buf_i2 = new_n963_;
  assign n519_i2 = ~new_n964_;
  assign n1029_i2 = new_n602_;
  assign n1041_i2 = new_n975_;
  assign n1043_i2 = new_n976_;
  assign n1045_i2 = new_n974_;
  assign n558_i2 = ~new_n977_;
  assign n563_i2 = ~new_n978_;
  assign lo094_buf_i2 = new_n616_;
  assign lo102_buf_i2 = new_n973_;
  assign n522_i2 = ~new_n979_;
  assign n527_i2 = ~new_n980_;
  assign n486_i2 = new_n981_;
  assign n491_i2 = new_n982_;
  assign n564_i2 = ~new_n757_;
  assign n528_i2 = ~new_n986_;
  assign n492_i2 = new_n994_;
  assign n530_i2 = ~new_n760_;
  assign n548_i2 = ~new_n761_;
  assign n536_i2 = ~new_n762_;
  assign n539_i2 = ~new_n763_;
  assign lo025_buf_i2 = new_n390_;
  assign lo073_buf_i2 = new_n420_;
  assign lo089_buf_i2 = new_n430_;
  assign lo121_buf_i2 = new_n452_;
  assign n509_i2 = new_n764_;
  assign n513_i2 = ~new_n766_;
  assign n501_i2 = ~new_n768_;
  assign n504_i2 = ~new_n770_;
  assign n495_i2 = ~new_n772_;
  assign n497_i2 = new_n773_;
  assign n515_i2 = new_n774_;
  assign n506_i2 = new_n775_;
  assign lo010_buf_i2 = new_n380_;
  assign lo042_buf_i2 = new_n400_;
  assign lo058_buf_i2 = new_n410_;
  assign lo138_buf_i2 = new_n462_;
  assign lo014_buf_i2 = new_n314_;
  assign lo022_buf_i2 = new_n995_;
  assign lo030_buf_i2 = new_n322_;
  assign lo038_buf_i2 = new_n996_;
  assign lo046_buf_i2 = new_n330_;
  assign lo054_buf_i2 = new_n997_;
  assign lo126_buf_i2 = new_n370_;
  assign lo134_buf_i2 = new_n998_;
  assign lo093_buf_i2 = new_n354_;
  assign lo101_buf_i2 = new_n358_;
  assign lo002_buf_i2 = new_n308_;
  assign lo006_buf_i2 = new_n310_;
  assign lo062_buf_i2 = new_n338_;
  assign lo070_buf_i2 = new_n342_;
  assign lo078_buf_i2 = new_n346_;
  assign lo086_buf_i2 = new_n350_;
  assign lo110_buf_i2 = new_n362_;
  assign lo118_buf_i2 = new_n366_;
  assign n476_i2 = new_n776_;
  assign n482_i2 = new_n777_;
  assign n478_i2 = new_n778_;
  assign n479_i2 = new_n779_;
  assign new_n919_ = new_n555_;
  assign new_n920_ = new_n919_;
  assign new_n921_ = new_n920_;
  assign new_n922_ = new_n919_;
  assign new_n923_ = new_n554_;
  assign new_n924_ = new_n923_;
  assign new_n925_ = new_n924_;
  assign new_n926_ = new_n924_;
  assign new_n927_ = new_n923_;
  assign new_n928_ = new_n927_;
  assign new_n929_ = new_n927_;
  assign new_n930_ = new_n650_;
  assign new_n931_ = new_n654_;
  assign new_n932_ = new_n657_;
  assign new_n933_ = new_n665_;
  assign new_n934_ = new_n664_;
  assign new_n935_ = new_n668_;
  assign new_n936_ = new_n673_;
  assign new_n937_ = new_n677_;
  assign new_n938_ = new_n679_;
  assign new_n939_ = new_n676_;
  assign new_n940_ = new_n684_;
  assign new_n941_ = new_n556_;
  assign new_n942_ = new_n941_;
  assign new_n943_ = new_n942_;
  assign new_n944_ = new_n941_;
  assign new_n945_ = new_n448_;
  assign new_n946_ = new_n706_;
  assign new_n947_ = new_n458_;
  assign new_n948_ = new_n704_;
  assign new_n949_ = new_n396_;
  assign new_n950_ = new_n698_;
  assign new_n951_ = new_n426_;
  assign new_n952_ = new_n700_;
  assign new_n953_ = new_n436_;
  assign new_n954_ = new_n702_;
  assign new_n955_ = new_n386_;
  assign new_n956_ = new_n693_;
  assign new_n957_ = new_n468_;
  assign new_n958_ = new_n696_;
  assign new_n959_ = new_n416_;
  assign new_n960_ = new_n695_;
  assign new_n961_ = new_n406_;
  assign new_n962_ = new_n694_;
  assign new_n963_ = new_n442_;
  assign new_n964_ = new_n712_;
  assign new_n965_ = new_n574_;
  assign new_n966_ = new_n710_;
  assign new_n967_ = new_n568_;
  assign new_n968_ = new_n707_;
  assign new_n969_ = new_n570_;
  assign new_n970_ = new_n708_;
  assign new_n971_ = new_n572_;
  assign new_n972_ = new_n709_;
  assign new_n973_ = new_n618_;
  assign new_n974_ = new_n634_;
  assign new_n975_ = new_n626_;
  assign new_n976_ = new_n630_;
  assign new_n977_ = new_n717_;
  assign new_n978_ = new_n728_;
  assign new_n979_ = new_n733_;
  assign new_n980_ = new_n744_;
  assign new_n981_ = new_n749_;
  assign new_n982_ = new_n756_;
  assign new_n983_ = new_n758_;
  assign new_n984_ = new_n983_;
  assign new_n985_ = new_n984_;
  assign new_n986_ = new_n983_;
  assign new_n987_ = new_n759_;
  assign new_n988_ = new_n987_;
  assign new_n989_ = new_n988_;
  assign new_n990_ = new_n989_;
  assign new_n991_ = new_n988_;
  assign new_n992_ = new_n987_;
  assign new_n993_ = new_n992_;
  assign new_n994_ = new_n992_;
  assign new_n995_ = new_n318_;
  assign new_n996_ = new_n326_;
  assign new_n997_ = new_n334_;
  assign new_n998_ = new_n374_;
  always @ (posedge clock) begin
    n229_lo <= n856_li008_li008;
    n253_lo <= n880_li016_li016;
    n256_lo <= n883_li017_li017;
    n259_lo <= n886_li018_li018;
    n262_lo <= n889_li019_li019;
    n277_lo <= n904_li024_li024;
    n301_lo <= n928_li032_li032;
    n304_lo <= n931_li033_li033;
    n307_lo <= n934_li034_li034;
    n310_lo <= n937_li035_li035;
    n325_lo <= n952_li040_li040;
    n349_lo <= n976_li048_li048;
    n352_lo <= n979_li049_li049;
    n355_lo <= n982_li050_li050;
    n358_lo <= n985_li051_li051;
    n373_lo <= n1000_li056_li056;
    n397_lo <= n1024_li064_li064;
    n400_lo <= n1027_li065_li065;
    n403_lo <= n1030_li066_li066;
    n406_lo <= n1033_li067_li067;
    n421_lo <= n1048_li072_li072;
    n445_lo <= n1072_li080_li080;
    n448_lo <= n1075_li081_li081;
    n451_lo <= n1078_li082_li082;
    n454_lo <= n1081_li083_li083;
    n469_lo <= n1096_li088_li088;
    n493_lo <= n1120_li096_li096;
    n496_lo <= n1123_li097_li097;
    n499_lo <= n1126_li098_li098;
    n502_lo <= n1129_li099_li099;
    n517_lo <= n1144_li104_li104;
    n520_lo <= n1147_li105_li105;
    n541_lo <= n1168_li112_li112;
    n544_lo <= n1171_li113_li113;
    n547_lo <= n1174_li114_li114;
    n550_lo <= n1177_li115_li115;
    n565_lo <= n1192_li120_li120;
    n589_lo <= n1216_li128_li128;
    n592_lo <= n1219_li129_li129;
    n595_lo <= n1222_li130_li130;
    n598_lo <= n1225_li131_li131;
    n613_lo <= n1240_li136_li136;
    n625_lo <= n1252_li140_li140;
    n628_lo <= n1255_li141_li141;
    n631_lo <= n1258_li142_li142;
    n634_lo <= n1261_li143_li143;
    n852_o2 <= n852_i2;
    n853_o2 <= n853_i2;
    n955_o2 <= n955_i2;
    n956_o2 <= n956_i2;
    n531_o2 <= n531_i2;
    n549_o2 <= n549_i2;
    n537_o2 <= n537_i2;
    n540_o2 <= n540_i2;
    n546_o2 <= n546_i2;
    n534_o2 <= n534_i2;
    n552_o2 <= n552_i2;
    n543_o2 <= n543_i2;
    n961_o2 <= n961_i2;
    n223_inv <= n962_i2;
    n555_o2 <= n555_i2;
    n1009_o2 <= n1009_i2;
    n1010_o2 <= n1010_i2;
    n1011_o2 <= n1011_i2;
    n1012_o2 <= n1012_i2;
    lo026_buf_o2 <= lo026_buf_i2;
    lo074_buf_o2 <= lo074_buf_i2;
    lo090_buf_o2 <= lo090_buf_i2;
    lo122_buf_o2 <= lo122_buf_i2;
    n510_o2 <= n510_i2;
    n498_o2 <= n498_i2;
    n516_o2 <= n516_i2;
    n507_o2 <= n507_i2;
    lo106_buf_o2 <= lo106_buf_i2;
    n519_o2 <= n519_i2;
    n1029_o2 <= n1029_i2;
    n1041_o2 <= n1041_i2;
    n1043_o2 <= n1043_i2;
    n1045_o2 <= n1045_i2;
    n558_o2 <= n558_i2;
    n563_o2 <= n563_i2;
    lo094_buf_o2 <= lo094_buf_i2;
    lo102_buf_o2 <= lo102_buf_i2;
    n522_o2 <= n522_i2;
    n298_inv <= n527_i2;
    n486_o2 <= n486_i2;
    n304_inv <= n491_i2;
    n564_o2 <= n564_i2;
    n528_o2 <= n528_i2;
    n492_o2 <= n492_i2;
    n530_o2 <= n530_i2;
    n548_o2 <= n548_i2;
    n536_o2 <= n536_i2;
    n539_o2 <= n539_i2;
    lo025_buf_o2 <= lo025_buf_i2;
    lo073_buf_o2 <= lo073_buf_i2;
    lo089_buf_o2 <= lo089_buf_i2;
    lo121_buf_o2 <= lo121_buf_i2;
    n509_o2 <= n509_i2;
    n513_o2 <= n513_i2;
    n501_o2 <= n501_i2;
    n504_o2 <= n504_i2;
    n495_o2 <= n495_i2;
    n497_o2 <= n497_i2;
    n515_o2 <= n515_i2;
    n506_o2 <= n506_i2;
    lo010_buf_o2 <= lo010_buf_i2;
    lo042_buf_o2 <= lo042_buf_i2;
    lo058_buf_o2 <= lo058_buf_i2;
    lo138_buf_o2 <= lo138_buf_i2;
    lo014_buf_o2 <= lo014_buf_i2;
    lo022_buf_o2 <= lo022_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo038_buf_o2 <= lo038_buf_i2;
    lo046_buf_o2 <= lo046_buf_i2;
    lo054_buf_o2 <= lo054_buf_i2;
    lo126_buf_o2 <= lo126_buf_i2;
    lo134_buf_o2 <= lo134_buf_i2;
    lo093_buf_o2 <= lo093_buf_i2;
    lo101_buf_o2 <= lo101_buf_i2;
    lo002_buf_o2 <= lo002_buf_i2;
    lo006_buf_o2 <= lo006_buf_i2;
    lo062_buf_o2 <= lo062_buf_i2;
    lo070_buf_o2 <= lo070_buf_i2;
    lo078_buf_o2 <= lo078_buf_i2;
    lo086_buf_o2 <= lo086_buf_i2;
    lo110_buf_o2 <= lo110_buf_i2;
    lo118_buf_o2 <= lo118_buf_i2;
    n476_o2 <= n476_i2;
    n482_o2 <= n482_i2;
    n478_o2 <= n478_i2;
    n479_o2 <= n479_i2;
  end
  initial begin
    n229_lo <= 1'b0;
    n253_lo <= 1'b0;
    n256_lo <= 1'b0;
    n259_lo <= 1'b0;
    n262_lo <= 1'b0;
    n277_lo <= 1'b0;
    n301_lo <= 1'b0;
    n304_lo <= 1'b0;
    n307_lo <= 1'b0;
    n310_lo <= 1'b0;
    n325_lo <= 1'b0;
    n349_lo <= 1'b0;
    n352_lo <= 1'b0;
    n355_lo <= 1'b0;
    n358_lo <= 1'b0;
    n373_lo <= 1'b0;
    n397_lo <= 1'b0;
    n400_lo <= 1'b0;
    n403_lo <= 1'b0;
    n406_lo <= 1'b0;
    n421_lo <= 1'b0;
    n445_lo <= 1'b0;
    n448_lo <= 1'b0;
    n451_lo <= 1'b0;
    n454_lo <= 1'b0;
    n469_lo <= 1'b0;
    n493_lo <= 1'b0;
    n496_lo <= 1'b0;
    n499_lo <= 1'b0;
    n502_lo <= 1'b0;
    n517_lo <= 1'b0;
    n520_lo <= 1'b0;
    n541_lo <= 1'b0;
    n544_lo <= 1'b0;
    n547_lo <= 1'b0;
    n550_lo <= 1'b0;
    n565_lo <= 1'b0;
    n589_lo <= 1'b0;
    n592_lo <= 1'b0;
    n595_lo <= 1'b0;
    n598_lo <= 1'b0;
    n613_lo <= 1'b0;
    n625_lo <= 1'b0;
    n628_lo <= 1'b0;
    n631_lo <= 1'b0;
    n634_lo <= 1'b0;
    n852_o2 <= 1'b0;
    n853_o2 <= 1'b0;
    n955_o2 <= 1'b0;
    n956_o2 <= 1'b0;
    n531_o2 <= 1'b0;
    n549_o2 <= 1'b0;
    n537_o2 <= 1'b0;
    n540_o2 <= 1'b0;
    n546_o2 <= 1'b0;
    n534_o2 <= 1'b0;
    n552_o2 <= 1'b0;
    n543_o2 <= 1'b0;
    n961_o2 <= 1'b0;
    n223_inv <= 1'b0;
    n555_o2 <= 1'b0;
    n1009_o2 <= 1'b0;
    n1010_o2 <= 1'b0;
    n1011_o2 <= 1'b0;
    n1012_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    n510_o2 <= 1'b0;
    n498_o2 <= 1'b0;
    n516_o2 <= 1'b0;
    n507_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n519_o2 <= 1'b0;
    n1029_o2 <= 1'b0;
    n1041_o2 <= 1'b0;
    n1043_o2 <= 1'b0;
    n1045_o2 <= 1'b0;
    n558_o2 <= 1'b0;
    n563_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    n522_o2 <= 1'b0;
    n298_inv <= 1'b0;
    n486_o2 <= 1'b0;
    n304_inv <= 1'b0;
    n564_o2 <= 1'b0;
    n528_o2 <= 1'b0;
    n492_o2 <= 1'b0;
    n530_o2 <= 1'b0;
    n548_o2 <= 1'b0;
    n536_o2 <= 1'b0;
    n539_o2 <= 1'b0;
    lo025_buf_o2 <= 1'b0;
    lo073_buf_o2 <= 1'b0;
    lo089_buf_o2 <= 1'b0;
    lo121_buf_o2 <= 1'b0;
    n509_o2 <= 1'b0;
    n513_o2 <= 1'b0;
    n501_o2 <= 1'b0;
    n504_o2 <= 1'b0;
    n495_o2 <= 1'b0;
    n497_o2 <= 1'b0;
    n515_o2 <= 1'b0;
    n506_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo138_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    lo134_buf_o2 <= 1'b0;
    lo093_buf_o2 <= 1'b0;
    lo101_buf_o2 <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    n476_o2 <= 1'b0;
    n482_o2 <= 1'b0;
    n478_o2 <= 1'b0;
    n479_o2 <= 1'b0;
  end
endmodule


